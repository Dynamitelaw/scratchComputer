module core ( gnd, vdd, clk, reset, instructionIn, start, busy, tempRegOut);

input gnd, vdd;
input clk;
input reset;
input start;
output busy;
input [31:0] instructionIn;
output [31:0] tempRegOut;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf9) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf8) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf7) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
	BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
	BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
	BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf8) );
	BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf7) );
	BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf6) );
	BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf5) );
	BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf4) );
	BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf3) );
	BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf2) );
	BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf1) );
	BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(_19153_), .Y(_19153__hier0_bF_buf0) );
	BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_20622_), .Y(_20622__bF_buf4) );
	BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(_20622_), .Y(_20622__bF_buf3) );
	BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(_20622_), .Y(_20622__bF_buf2) );
	BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(_20622_), .Y(_20622__bF_buf1) );
	BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(_20622_), .Y(_20622__bF_buf0) );
	BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(_17412_), .Y(_17412__bF_buf4) );
	BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(_17412_), .Y(_17412__bF_buf3) );
	BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_17412_), .Y(_17412__bF_buf2) );
	BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_17412_), .Y(_17412__bF_buf1) );
	BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_17412_), .Y(_17412__bF_buf0) );
	BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_20580_), .Y(_20580__bF_buf4) );
	BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_20580_), .Y(_20580__bF_buf3) );
	BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_20580_), .Y(_20580__bF_buf2) );
	BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_20580_), .Y(_20580__bF_buf1) );
	BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_20580_), .Y(_20580__bF_buf0) );
	BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_), .Y(reg_dataIn_31_bF_buf4) );
	BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_), .Y(reg_dataIn_31_bF_buf3) );
	BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_), .Y(reg_dataIn_31_bF_buf2) );
	BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_), .Y(reg_dataIn_31_bF_buf1) );
	BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_), .Y(reg_dataIn_31_bF_buf0) );
	BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract), .Y(adder_subtract_bF_buf3) );
	BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract), .Y(adder_subtract_bF_buf2) );
	BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract), .Y(adder_subtract_bF_buf1) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract), .Y(adder_subtract_bF_buf0) );
	BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .Y(_3263__bF_buf3) );
	BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .Y(_3263__bF_buf2) );
	BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .Y(_3263__bF_buf1) );
	BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .Y(_3263__bF_buf0) );
	BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_), .Y(divider_absoluteValue_B_flipSign_result_26_bF_buf3) );
	BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_), .Y(divider_absoluteValue_B_flipSign_result_26_bF_buf2) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_), .Y(divider_absoluteValue_B_flipSign_result_26_bF_buf1) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_), .Y(divider_absoluteValue_B_flipSign_result_26_bF_buf0) );
	BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[31]), .Y(instructionIn_31_bF_buf3) );
	BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[31]), .Y(instructionIn_31_bF_buf2) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[31]), .Y(instructionIn_31_bF_buf1) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[31]), .Y(instructionIn_31_bF_buf0) );
	BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf7) );
	BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf6) );
	BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf5) );
	BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf4) );
	BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf3) );
	BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf2) );
	BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf1) );
	BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_19292_), .Y(_19292__bF_buf0) );
	BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_), .Y(aOperand_frameOut_16_bF_buf4) );
	BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_), .Y(aOperand_frameOut_16_bF_buf3) );
	BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_), .Y(aOperand_frameOut_16_bF_buf2) );
	BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_), .Y(aOperand_frameOut_16_bF_buf1) );
	BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_), .Y(aOperand_frameOut_16_bF_buf0) );
	BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf7) );
	BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf6) );
	BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf5) );
	BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf4) );
	BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf3) );
	BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf2) );
	BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf1) );
	BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_19533_), .Y(_19533__bF_buf0) );
	BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .Y(_12310__bF_buf3) );
	BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .Y(_12310__bF_buf2) );
	BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .Y(_12310__bF_buf1) );
	BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .Y(_12310__bF_buf0) );
	BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf7) );
	BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf6) );
	BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf5) );
	BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf4) );
	BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf3) );
	BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf2) );
	BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf1) );
	BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(_19804_), .Y(_19804__bF_buf0) );
	BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(_17236_), .Y(_17236__bF_buf3) );
	BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(_17236_), .Y(_17236__bF_buf2) );
	BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(_17236_), .Y(_17236__bF_buf1) );
	BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(_17236_), .Y(_17236__bF_buf0) );
	BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_), .Y(reg_dataIn_29_bF_buf4) );
	BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_), .Y(reg_dataIn_29_bF_buf3) );
	BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_), .Y(reg_dataIn_29_bF_buf2) );
	BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_), .Y(reg_dataIn_29_bF_buf1) );
	BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_), .Y(reg_dataIn_29_bF_buf0) );
	BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(_20615_), .Y(_20615__bF_buf4) );
	BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(_20615_), .Y(_20615__bF_buf3) );
	BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_20615_), .Y(_20615__bF_buf2) );
	BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_20615_), .Y(_20615__bF_buf1) );
	BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(_20615_), .Y(_20615__bF_buf0) );
	BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf7) );
	BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf6) );
	BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf5) );
	BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf4) );
	BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf3) );
	BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf2) );
	BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf1) );
	BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(_19702_), .Y(_19702__bF_buf0) );
	BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_17435_), .Y(_17435__bF_buf4) );
	BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_17435_), .Y(_17435__bF_buf3) );
	BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_17435_), .Y(_17435__bF_buf2) );
	BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_17435_), .Y(_17435__bF_buf1) );
	BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(_17435_), .Y(_17435__bF_buf0) );
	BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf6) );
	BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf5) );
	BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf4) );
	BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf3) );
	BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf2) );
	BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf1) );
	BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_8052_), .Y(_8052__bF_buf0) );
	BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_), .Y(divider_absoluteValue_B_flipSign_result_21_bF_buf3) );
	BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_), .Y(divider_absoluteValue_B_flipSign_result_21_bF_buf2) );
	BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_), .Y(divider_absoluteValue_B_flipSign_result_21_bF_buf1) );
	BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_), .Y(divider_absoluteValue_B_flipSign_result_21_bF_buf0) );
	BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(_17393_), .Y(_17393__bF_buf4) );
	BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(_17393_), .Y(_17393__bF_buf3) );
	BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(_17393_), .Y(_17393__bF_buf2) );
	BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(_17393_), .Y(_17393__bF_buf1) );
	BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(_17393_), .Y(_17393__bF_buf0) );
	BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_), .Y(aOperand_frameOut_11_bF_buf4) );
	BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_), .Y(aOperand_frameOut_11_bF_buf3) );
	BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_), .Y(aOperand_frameOut_11_bF_buf2) );
	BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_), .Y(aOperand_frameOut_11_bF_buf1) );
	BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_), .Y(aOperand_frameOut_11_bF_buf0) );
	BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_), .Y(aOperand_frameOut_6_bF_buf4) );
	BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_), .Y(aOperand_frameOut_6_bF_buf3) );
	BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_), .Y(aOperand_frameOut_6_bF_buf2) );
	BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_), .Y(aOperand_frameOut_6_bF_buf1) );
	BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_), .Y(aOperand_frameOut_6_bF_buf0) );
	BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_), .Y(reg_dataIn_24_bF_buf4) );
	BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_), .Y(reg_dataIn_24_bF_buf3) );
	BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_), .Y(reg_dataIn_24_bF_buf2) );
	BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_), .Y(reg_dataIn_24_bF_buf1) );
	BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_), .Y(reg_dataIn_24_bF_buf0) );
	BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_20610_), .Y(_20610__bF_buf4) );
	BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(_20610_), .Y(_20610__bF_buf3) );
	BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(_20610_), .Y(_20610__bF_buf2) );
	BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(_20610_), .Y(_20610__bF_buf1) );
	BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(_20610_), .Y(_20610__bF_buf0) );
	BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(_17400_), .Y(_17400__bF_buf4) );
	BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(_17400_), .Y(_17400__bF_buf3) );
	BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(_17400_), .Y(_17400__bF_buf2) );
	BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(_17400_), .Y(_17400__bF_buf1) );
	BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(_17400_), .Y(_17400__bF_buf0) );
	BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf106) );
	BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf105) );
	BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf104) );
	BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf103) );
	BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf102) );
	BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf101) );
	BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf100) );
	BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf99) );
	BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf98) );
	BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf97) );
	BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf96) );
	BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf95) );
	BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf94) );
	BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf93) );
	BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf92) );
	BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf91) );
	BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf90) );
	BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf89) );
	BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf88) );
	BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf87) );
	BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf86) );
	BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf85) );
	BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf84) );
	BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf83) );
	BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf82) );
	BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf81) );
	BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf80) );
	BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf79) );
	BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf78) );
	BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf77) );
	BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf76) );
	BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf75) );
	BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf74) );
	BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf73) );
	BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf72) );
	BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf71) );
	BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf70) );
	BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf69) );
	BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf68) );
	BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf67) );
	BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf66) );
	BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf65) );
	BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf64) );
	BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf63) );
	BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf62) );
	BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf61) );
	BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf60) );
	BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf59) );
	BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf58) );
	BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf57) );
	BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf56) );
	BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf55) );
	BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf54) );
	BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf53) );
	BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf52) );
	BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf51) );
	BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf50) );
	BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf49) );
	BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf48) );
	BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf47) );
	BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf46) );
	BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf45) );
	BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf44) );
	BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf43) );
	BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf42) );
	BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf41) );
	BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf40) );
	BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf39) );
	BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf38) );
	BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf37) );
	BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf36) );
	BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf35) );
	BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf34) );
	BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf33) );
	BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf32) );
	BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf31) );
	BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf30) );
	BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf29) );
	BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28) );
	BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf27) );
	BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf26) );
	BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf25) );
	BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf24) );
	BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf23) );
	BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf22) );
	BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf21) );
	BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf20) );
	BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf19) );
	BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf18) );
	BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf17) );
	BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf16) );
	BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf15) );
	BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf14) );
	BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf13) );
	BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf12) );
	BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_), .Y(aOperand_frameOut_1_bF_buf5) );
	BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_), .Y(aOperand_frameOut_1_bF_buf4) );
	BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_), .Y(aOperand_frameOut_1_bF_buf3) );
	BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_), .Y(aOperand_frameOut_1_bF_buf2) );
	BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_), .Y(aOperand_frameOut_1_bF_buf1) );
	BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_), .Y(aOperand_frameOut_1_bF_buf0) );
	BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .Y(_13294__bF_buf3) );
	BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .Y(_13294__bF_buf2) );
	BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .Y(_13294__bF_buf1) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_13294_), .Y(_13294__bF_buf0) );
	BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_), .Y(divider_absoluteValue_B_flipSign_result_19_bF_buf4) );
	BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_), .Y(divider_absoluteValue_B_flipSign_result_19_bF_buf3) );
	BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_), .Y(divider_absoluteValue_B_flipSign_result_19_bF_buf2) );
	BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_), .Y(divider_absoluteValue_B_flipSign_result_19_bF_buf1) );
	BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_), .Y(divider_absoluteValue_B_flipSign_result_19_bF_buf0) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_), .Y(adder_bOperand_17_bF_buf3) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_), .Y(adder_bOperand_17_bF_buf2) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_), .Y(adder_bOperand_17_bF_buf1) );
	BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_), .Y(adder_bOperand_17_bF_buf0) );
	BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf3) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf2) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf1) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_4881_), .Y(_4881__bF_buf0) );
	BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .Y(_11636__bF_buf4) );
	BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .Y(_11636__bF_buf3) );
	BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .Y(_11636__bF_buf2) );
	BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .Y(_11636__bF_buf1) );
	BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(_11636_), .Y(_11636__bF_buf0) );
	BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_), .Y(reg_dataIn_7_bF_buf4) );
	BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_), .Y(reg_dataIn_7_bF_buf3) );
	BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_), .Y(reg_dataIn_7_bF_buf2) );
	BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_), .Y(reg_dataIn_7_bF_buf1) );
	BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_), .Y(reg_dataIn_7_bF_buf0) );
	BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf7) );
	BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf6) );
	BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf5) );
	BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf4) );
	BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf3) );
	BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf2) );
	BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf1) );
	BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(_20066_), .Y(_20066__bF_buf0) );
	BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf98) );
	BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf97) );
	BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf96) );
	BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf95) );
	BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf94) );
	BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf93) );
	BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf92) );
	BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf91) );
	BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf90) );
	BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf89) );
	BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf88) );
	BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf87) );
	BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf86) );
	BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf85) );
	BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf84) );
	BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf83) );
	BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf82) );
	BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf81) );
	BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf80) );
	BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf79) );
	BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf78) );
	BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf77) );
	BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf76) );
	BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf75) );
	BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf74) );
	BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf73) );
	BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf72) );
	BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf71) );
	BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf70) );
	BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf69) );
	BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf68) );
	BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf67) );
	BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf66) );
	BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf65) );
	BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf64) );
	BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf63) );
	BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf62) );
	BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf61) );
	BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf60) );
	BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf59) );
	BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf58) );
	BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf57) );
	BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf56) );
	BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf55) );
	BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf54) );
	BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf53) );
	BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf52) );
	BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf51) );
	BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf50) );
	BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf49) );
	BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf48) );
	BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf47) );
	BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf46) );
	BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf45) );
	BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf44) );
	BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf43) );
	BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf42) );
	BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf41) );
	BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf40) );
	BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf39) );
	BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf38) );
	BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf37) );
	BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf36) );
	BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf35) );
	BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf34) );
	BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf33) );
	BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf32) );
	BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf31) );
	BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf30) );
	BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf29) );
	BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf28) );
	BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf27) );
	BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf26) );
	BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf25) );
	BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf24) );
	BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf23) );
	BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf22) );
	BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf21) );
	BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf20) );
	BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf19) );
	BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf18) );
	BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf17) );
	BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf16) );
	BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf15) );
	BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf14) );
	BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf13) );
	BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf12) );
	BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf11) );
	BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf10) );
	BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf9) );
	BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf8), .Y(_19153__bF_buf8) );
	BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf7), .Y(_19153__bF_buf7) );
	BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf6), .Y(_19153__bF_buf6) );
	BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf5), .Y(_19153__bF_buf5) );
	BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf4), .Y(_19153__bF_buf4) );
	BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf3), .Y(_19153__bF_buf3) );
	BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf2), .Y(_19153__bF_buf2) );
	BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf1), .Y(_19153__bF_buf1) );
	BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(_19153__hier0_bF_buf0), .Y(_19153__bF_buf0) );
	BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1484__bF_buf4) );
	BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1484__bF_buf3) );
	BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1484__bF_buf2) );
	BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1484__bF_buf1) );
	BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .Y(_1484__bF_buf0) );
	BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(_20608_), .Y(_20608__bF_buf4) );
	BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(_20608_), .Y(_20608__bF_buf3) );
	BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(_20608_), .Y(_20608__bF_buf2) );
	BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(_20608_), .Y(_20608__bF_buf1) );
	BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(_20608_), .Y(_20608__bF_buf0) );
	BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_78__bF_buf4) );
	BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_78__bF_buf3) );
	BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_78__bF_buf2) );
	BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_78__bF_buf1) );
	BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_78__bF_buf0) );
	BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_), .Y(divider_absoluteValue_B_flipSign_result_14_bF_buf5) );
	BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_), .Y(divider_absoluteValue_B_flipSign_result_14_bF_buf4) );
	BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_), .Y(divider_absoluteValue_B_flipSign_result_14_bF_buf3) );
	BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_), .Y(divider_absoluteValue_B_flipSign_result_14_bF_buf2) );
	BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_), .Y(divider_absoluteValue_B_flipSign_result_14_bF_buf1) );
	BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_), .Y(divider_absoluteValue_B_flipSign_result_14_bF_buf0) );
	BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .Y(_2922__bF_buf3) );
	BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .Y(_2922__bF_buf2) );
	BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .Y(_2922__bF_buf1) );
	BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .Y(_2922__bF_buf0) );
	BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_), .Y(adder_bOperand_12_bF_buf3) );
	BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_), .Y(adder_bOperand_12_bF_buf2) );
	BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_), .Y(adder_bOperand_12_bF_buf1) );
	BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_), .Y(adder_bOperand_12_bF_buf0) );
	BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(_17025_), .Y(_17025__bF_buf3) );
	BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(_17025_), .Y(_17025__bF_buf2) );
	BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(_17025_), .Y(_17025__bF_buf1) );
	BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(_17025_), .Y(_17025__bF_buf0) );
	BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf7) );
	BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf6) );
	BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf5) );
	BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf4) );
	BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf3) );
	BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf2) );
	BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf1) );
	BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(_19220_), .Y(_19220__bF_buf0) );
	BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_), .Y(reg_dataIn_2_bF_buf4) );
	BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_), .Y(reg_dataIn_2_bF_buf3) );
	BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_), .Y(reg_dataIn_2_bF_buf2) );
	BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_), .Y(reg_dataIn_2_bF_buf1) );
	BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_), .Y(reg_dataIn_2_bF_buf0) );
	BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_), .Y(reg_dataIn_17_bF_buf4) );
	BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_), .Y(reg_dataIn_17_bF_buf3) );
	BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_), .Y(reg_dataIn_17_bF_buf2) );
	BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_), .Y(reg_dataIn_17_bF_buf1) );
	BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_), .Y(reg_dataIn_17_bF_buf0) );
	BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf8) );
	BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf7) );
	BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf6) );
	BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf5) );
	BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf4) );
	BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf3) );
	BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf2) );
	BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf1) );
	BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative), .Y(divider_a_isNegative_bF_buf0) );
	BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(_20633_), .Y(_20633__bF_buf4) );
	BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(_20633_), .Y(_20633__bF_buf3) );
	BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(_20633_), .Y(_20633__bF_buf2) );
	BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(_20633_), .Y(_20633__bF_buf1) );
	BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(_20633_), .Y(_20633__bF_buf0) );
	BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf6) );
	BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf5) );
	BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf4) );
	BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf3) );
	BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf2) );
	BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf1) );
	BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_), .Y(divider_absoluteValue_B_flipSign_result_7_bF_buf0) );
	BUFX4 BUFX4_464 ( .gnd(gnd), .vdd(vdd), .A(_17423_), .Y(_17423__bF_buf4) );
	BUFX4 BUFX4_465 ( .gnd(gnd), .vdd(vdd), .A(_17423_), .Y(_17423__bF_buf3) );
	BUFX4 BUFX4_466 ( .gnd(gnd), .vdd(vdd), .A(_17423_), .Y(_17423__bF_buf2) );
	BUFX4 BUFX4_467 ( .gnd(gnd), .vdd(vdd), .A(_17423_), .Y(_17423__bF_buf1) );
	BUFX4 BUFX4_468 ( .gnd(gnd), .vdd(vdd), .A(_17423_), .Y(_17423__bF_buf0) );
	BUFX4 BUFX4_469 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .Y(_5377__bF_buf5) );
	BUFX4 BUFX4_470 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .Y(_5377__bF_buf4) );
	BUFX4 BUFX4_471 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .Y(_5377__bF_buf3) );
	BUFX4 BUFX4_472 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .Y(_5377__bF_buf2) );
	BUFX4 BUFX4_473 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .Y(_5377__bF_buf1) );
	BUFX4 BUFX4_474 ( .gnd(gnd), .vdd(vdd), .A(_5377_), .Y(_5377__bF_buf0) );
	BUFX4 BUFX4_475 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .Y(_6315__bF_buf5) );
	BUFX4 BUFX4_476 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .Y(_6315__bF_buf4) );
	BUFX4 BUFX4_477 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .Y(_6315__bF_buf3) );
	BUFX4 BUFX4_478 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .Y(_6315__bF_buf2) );
	BUFX4 BUFX4_479 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .Y(_6315__bF_buf1) );
	BUFX4 BUFX4_480 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .Y(_6315__bF_buf0) );
	BUFX4 BUFX4_481 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_), .Y(adder_bOperand_8_bF_buf4) );
	BUFX4 BUFX4_482 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_), .Y(adder_bOperand_8_bF_buf3) );
	BUFX4 BUFX4_483 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_), .Y(adder_bOperand_8_bF_buf2) );
	BUFX4 BUFX4_484 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_), .Y(adder_bOperand_8_bF_buf1) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_), .Y(adder_bOperand_8_bF_buf0) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_5516_), .Y(_5516__bF_buf3) );
	BUFX4 BUFX4_485 ( .gnd(gnd), .vdd(vdd), .A(_5516_), .Y(_5516__bF_buf2) );
	BUFX4 BUFX4_486 ( .gnd(gnd), .vdd(vdd), .A(_5516_), .Y(_5516__bF_buf1) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_5516_), .Y(_5516__bF_buf0) );
	BUFX4 BUFX4_487 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_), .Y(reg_dataIn_12_bF_buf4) );
	BUFX4 BUFX4_488 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_), .Y(reg_dataIn_12_bF_buf3) );
	BUFX4 BUFX4_489 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_), .Y(reg_dataIn_12_bF_buf2) );
	BUFX4 BUFX4_490 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_), .Y(reg_dataIn_12_bF_buf1) );
	BUFX4 BUFX4_491 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_), .Y(reg_dataIn_12_bF_buf0) );
	BUFX4 BUFX4_492 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_), .Y(divider_divuResult_15_bF_buf4) );
	BUFX4 BUFX4_493 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_), .Y(divider_divuResult_15_bF_buf3) );
	BUFX4 BUFX4_494 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_), .Y(divider_divuResult_15_bF_buf2) );
	BUFX4 BUFX4_495 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_), .Y(divider_divuResult_15_bF_buf1) );
	BUFX4 BUFX4_496 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_), .Y(divider_divuResult_15_bF_buf0) );
	BUFX4 BUFX4_497 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf7) );
	BUFX4 BUFX4_498 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf6) );
	BUFX4 BUFX4_499 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf5) );
	BUFX4 BUFX4_500 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf4) );
	BUFX4 BUFX4_501 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf3) );
	BUFX4 BUFX4_502 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf2) );
	BUFX4 BUFX4_503 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf1) );
	BUFX4 BUFX4_504 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_), .Y(divider_absoluteValue_B_flipSign_result_2_bF_buf0) );
	BUFX4 BUFX4_505 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_), .Y(adder_bOperand_3_bF_buf5) );
	BUFX4 BUFX4_506 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_), .Y(adder_bOperand_3_bF_buf4) );
	BUFX4 BUFX4_507 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_), .Y(adder_bOperand_3_bF_buf3) );
	BUFX4 BUFX4_508 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_), .Y(adder_bOperand_3_bF_buf2) );
	BUFX4 BUFX4_509 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_), .Y(adder_bOperand_3_bF_buf1) );
	BUFX4 BUFX4_510 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_), .Y(adder_bOperand_3_bF_buf0) );
	BUFX4 BUFX4_511 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf6) );
	BUFX4 BUFX4_512 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf5) );
	BUFX4 BUFX4_513 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf4) );
	BUFX4 BUFX4_514 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf3) );
	BUFX4 BUFX4_515 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf2) );
	BUFX4 BUFX4_516 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf1) );
	BUFX4 BUFX4_517 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .Y(_6840__bF_buf0) );
	BUFX4 BUFX4_518 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf7) );
	BUFX4 BUFX4_519 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf6) );
	BUFX4 BUFX4_520 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf5) );
	BUFX4 BUFX4_521 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf4) );
	BUFX4 BUFX4_522 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf3) );
	BUFX4 BUFX4_523 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf2) );
	BUFX4 BUFX4_524 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf1) );
	BUFX4 BUFX4_525 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .Y(_2547__bF_buf0) );
	BUFX4 BUFX4_526 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_), .Y(divider_divuResult_10_bF_buf5) );
	BUFX4 BUFX4_527 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_), .Y(divider_divuResult_10_bF_buf4) );
	BUFX4 BUFX4_528 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_), .Y(divider_divuResult_10_bF_buf3) );
	BUFX4 BUFX4_529 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_), .Y(divider_divuResult_10_bF_buf2) );
	BUFX4 BUFX4_530 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_), .Y(divider_divuResult_10_bF_buf1) );
	BUFX4 BUFX4_531 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_), .Y(divider_divuResult_10_bF_buf0) );
	BUFX4 BUFX4_532 ( .gnd(gnd), .vdd(vdd), .A(_20589_), .Y(_20589__bF_buf4) );
	BUFX4 BUFX4_533 ( .gnd(gnd), .vdd(vdd), .A(_20589_), .Y(_20589__bF_buf3) );
	BUFX4 BUFX4_534 ( .gnd(gnd), .vdd(vdd), .A(_20589_), .Y(_20589__bF_buf2) );
	BUFX4 BUFX4_535 ( .gnd(gnd), .vdd(vdd), .A(_20589_), .Y(_20589__bF_buf1) );
	BUFX4 BUFX4_536 ( .gnd(gnd), .vdd(vdd), .A(_20589_), .Y(_20589__bF_buf0) );
	BUFX4 BUFX4_537 ( .gnd(gnd), .vdd(vdd), .A(_20559_), .Y(_20559__bF_buf5) );
	BUFX4 BUFX4_538 ( .gnd(gnd), .vdd(vdd), .A(_20559_), .Y(_20559__bF_buf4) );
	BUFX4 BUFX4_539 ( .gnd(gnd), .vdd(vdd), .A(_20559_), .Y(_20559__bF_buf3) );
	BUFX4 BUFX4_540 ( .gnd(gnd), .vdd(vdd), .A(_20559_), .Y(_20559__bF_buf2) );
	BUFX4 BUFX4_541 ( .gnd(gnd), .vdd(vdd), .A(_20559_), .Y(_20559__bF_buf1) );
	BUFX4 BUFX4_542 ( .gnd(gnd), .vdd(vdd), .A(_20559_), .Y(_20559__bF_buf0) );
	BUFX4 BUFX4_543 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .Y(_2042__bF_buf3) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .Y(_2042__bF_buf2) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .Y(_2042__bF_buf1) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .Y(_2042__bF_buf0) );
	BUFX4 BUFX4_544 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf6) );
	BUFX4 BUFX4_545 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf5) );
	BUFX4 BUFX4_546 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf4) );
	BUFX4 BUFX4_547 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf3) );
	BUFX4 BUFX4_548 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf2) );
	BUFX4 BUFX4_549 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf1) );
	BUFX4 BUFX4_550 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_), .Y(divider_divuResult_6_bF_buf0) );
	BUFX4 BUFX4_551 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf7) );
	BUFX4 BUFX4_552 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf6) );
	BUFX4 BUFX4_553 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf5) );
	BUFX4 BUFX4_554 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf4) );
	BUFX4 BUFX4_555 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf3) );
	BUFX4 BUFX4_556 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf2) );
	BUFX4 BUFX4_557 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf1) );
	BUFX4 BUFX4_558 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .Y(_2470__bF_buf0) );
	BUFX4 BUFX4_559 ( .gnd(gnd), .vdd(vdd), .A(_20626_), .Y(_20626__bF_buf4) );
	BUFX4 BUFX4_560 ( .gnd(gnd), .vdd(vdd), .A(_20626_), .Y(_20626__bF_buf3) );
	BUFX4 BUFX4_561 ( .gnd(gnd), .vdd(vdd), .A(_20626_), .Y(_20626__bF_buf2) );
	BUFX4 BUFX4_562 ( .gnd(gnd), .vdd(vdd), .A(_20626_), .Y(_20626__bF_buf1) );
	BUFX4 BUFX4_563 ( .gnd(gnd), .vdd(vdd), .A(_20626_), .Y(_20626__bF_buf0) );
	BUFX4 BUFX4_564 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .Y(_10855__bF_buf4) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .Y(_10855__bF_buf3) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .Y(_10855__bF_buf2) );
	BUFX4 BUFX4_565 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .Y(_10855__bF_buf1) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_10855_), .Y(_10855__bF_buf0) );
	BUFX4 BUFX4_566 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_66__bF_buf4) );
	BUFX4 BUFX4_567 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_66__bF_buf3) );
	BUFX4 BUFX4_568 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_66__bF_buf2) );
	BUFX4 BUFX4_569 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_66__bF_buf1) );
	BUFX4 BUFX4_570 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_66__bF_buf0) );
	BUFX4 BUFX4_571 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .Y(_11450__bF_buf4) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .Y(_11450__bF_buf3) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .Y(_11450__bF_buf2) );
	BUFX4 BUFX4_572 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .Y(_11450__bF_buf1) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .Y(_11450__bF_buf0) );
	BUFX4 BUFX4_573 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf6) );
	BUFX4 BUFX4_574 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf5) );
	BUFX4 BUFX4_575 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf4) );
	BUFX4 BUFX4_576 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf3) );
	BUFX4 BUFX4_577 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf2) );
	BUFX4 BUFX4_578 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf1) );
	BUFX4 BUFX4_579 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_), .Y(divider_divuResult_1_bF_buf0) );
	BUFX4 BUFX4_580 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_), .Y(aOperand_frameOut_22_bF_buf3) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_), .Y(aOperand_frameOut_22_bF_buf2) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_), .Y(aOperand_frameOut_22_bF_buf1) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_), .Y(aOperand_frameOut_22_bF_buf0) );
	BUFX4 BUFX4_581 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf7) );
	BUFX4 BUFX4_582 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf6) );
	BUFX4 BUFX4_583 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf5) );
	BUFX4 BUFX4_584 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf4) );
	BUFX4 BUFX4_585 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf3) );
	BUFX4 BUFX4_586 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf2) );
	BUFX4 BUFX4_587 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf1) );
	BUFX4 BUFX4_588 ( .gnd(gnd), .vdd(vdd), .A(_19870_), .Y(_19870__bF_buf0) );
	BUFX4 BUFX4_589 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_7204__bF_buf5) );
	BUFX4 BUFX4_590 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_7204__bF_buf4) );
	BUFX4 BUFX4_591 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_7204__bF_buf3) );
	BUFX4 BUFX4_592 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_7204__bF_buf2) );
	BUFX4 BUFX4_593 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_7204__bF_buf1) );
	BUFX4 BUFX4_594 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_7204__bF_buf0) );
	BUFX4 BUFX4_595 ( .gnd(gnd), .vdd(vdd), .A(_20621_), .Y(_20621__bF_buf4) );
	BUFX4 BUFX4_596 ( .gnd(gnd), .vdd(vdd), .A(_20621_), .Y(_20621__bF_buf3) );
	BUFX4 BUFX4_597 ( .gnd(gnd), .vdd(vdd), .A(_20621_), .Y(_20621__bF_buf2) );
	BUFX4 BUFX4_598 ( .gnd(gnd), .vdd(vdd), .A(_20621_), .Y(_20621__bF_buf1) );
	BUFX4 BUFX4_599 ( .gnd(gnd), .vdd(vdd), .A(_20621_), .Y(_20621__bF_buf0) );
	BUFX4 BUFX4_600 ( .gnd(gnd), .vdd(vdd), .A(_17411_), .Y(_17411__bF_buf5) );
	BUFX4 BUFX4_601 ( .gnd(gnd), .vdd(vdd), .A(_17411_), .Y(_17411__bF_buf4) );
	BUFX4 BUFX4_602 ( .gnd(gnd), .vdd(vdd), .A(_17411_), .Y(_17411__bF_buf3) );
	BUFX4 BUFX4_603 ( .gnd(gnd), .vdd(vdd), .A(_17411_), .Y(_17411__bF_buf2) );
	BUFX4 BUFX4_604 ( .gnd(gnd), .vdd(vdd), .A(_17411_), .Y(_17411__bF_buf1) );
	BUFX4 BUFX4_605 ( .gnd(gnd), .vdd(vdd), .A(_17411_), .Y(_17411__bF_buf0) );
	BUFX4 BUFX4_606 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf6) );
	BUFX4 BUFX4_607 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf5) );
	BUFX4 BUFX4_608 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf4) );
	BUFX4 BUFX4_609 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf3) );
	BUFX4 BUFX4_610 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf2) );
	BUFX4 BUFX4_611 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf1) );
	BUFX4 BUFX4_612 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .Y(_4999__bF_buf0) );
	BUFX4 BUFX4_613 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_), .Y(reg_dataIn_30_bF_buf4) );
	BUFX4 BUFX4_614 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_), .Y(reg_dataIn_30_bF_buf3) );
	BUFX4 BUFX4_615 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_), .Y(reg_dataIn_30_bF_buf2) );
	BUFX4 BUFX4_616 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_), .Y(reg_dataIn_30_bF_buf1) );
	BUFX4 BUFX4_617 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_), .Y(reg_dataIn_30_bF_buf0) );
	BUFX4 BUFX4_618 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf4) );
	BUFX4 BUFX4_619 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf3) );
	BUFX4 BUFX4_620 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf2) );
	BUFX4 BUFX4_621 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf1) );
	BUFX4 BUFX4_622 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf0) );
	BUFX4 BUFX4_623 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf7) );
	BUFX4 BUFX4_624 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf6) );
	BUFX4 BUFX4_625 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf5) );
	BUFX4 BUFX4_626 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf4) );
	BUFX4 BUFX4_627 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf3) );
	BUFX4 BUFX4_628 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf2) );
	BUFX4 BUFX4_629 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf1) );
	BUFX4 BUFX4_630 ( .gnd(gnd), .vdd(vdd), .A(_19567_), .Y(_19567__bF_buf0) );
	BUFX4 BUFX4_631 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .Y(_3262__bF_buf4) );
	BUFX4 BUFX4_632 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .Y(_3262__bF_buf3) );
	BUFX4 BUFX4_633 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .Y(_3262__bF_buf2) );
	BUFX4 BUFX4_634 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .Y(_3262__bF_buf1) );
	BUFX4 BUFX4_635 ( .gnd(gnd), .vdd(vdd), .A(_3262_), .Y(_3262__bF_buf0) );
	BUFX4 BUFX4_636 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf7) );
	BUFX4 BUFX4_637 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf6) );
	BUFX4 BUFX4_638 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf5) );
	BUFX4 BUFX4_639 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf4) );
	BUFX4 BUFX4_640 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf3) );
	BUFX4 BUFX4_641 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf2) );
	BUFX4 BUFX4_642 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf1) );
	BUFX4 BUFX4_643 ( .gnd(gnd), .vdd(vdd), .A(_19736_), .Y(_19736__bF_buf0) );
	BUFX4 BUFX4_644 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf6) );
	BUFX4 BUFX4_645 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf5) );
	BUFX4 BUFX4_646 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf4) );
	BUFX4 BUFX4_647 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf3) );
	BUFX4 BUFX4_648 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf2) );
	BUFX4 BUFX4_649 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf1) );
	BUFX4 BUFX4_650 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9325__bF_buf0) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_), .Y(aOperand_frameOut_15_bF_buf4) );
	BUFX4 BUFX4_651 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_), .Y(aOperand_frameOut_15_bF_buf3) );
	BUFX4 BUFX4_652 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_), .Y(aOperand_frameOut_15_bF_buf2) );
	BUFX4 BUFX4_653 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_), .Y(aOperand_frameOut_15_bF_buf1) );
	BUFX4 BUFX4_654 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_), .Y(aOperand_frameOut_15_bF_buf0) );
	BUFX4 BUFX4_655 ( .gnd(gnd), .vdd(vdd), .A(_17295_), .Y(_17295__bF_buf4) );
	BUFX4 BUFX4_656 ( .gnd(gnd), .vdd(vdd), .A(_17295_), .Y(_17295__bF_buf3) );
	BUFX4 BUFX4_657 ( .gnd(gnd), .vdd(vdd), .A(_17295_), .Y(_17295__bF_buf2) );
	BUFX4 BUFX4_658 ( .gnd(gnd), .vdd(vdd), .A(_17295_), .Y(_17295__bF_buf1) );
	BUFX4 BUFX4_659 ( .gnd(gnd), .vdd(vdd), .A(_17295_), .Y(_17295__bF_buf0) );
	BUFX4 BUFX4_660 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_), .Y(reg_dataIn_28_bF_buf4) );
	BUFX4 BUFX4_661 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_), .Y(reg_dataIn_28_bF_buf3) );
	BUFX4 BUFX4_662 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_), .Y(reg_dataIn_28_bF_buf2) );
	BUFX4 BUFX4_663 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_), .Y(reg_dataIn_28_bF_buf1) );
	BUFX4 BUFX4_664 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_), .Y(reg_dataIn_28_bF_buf0) );
	BUFX4 BUFX4_665 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_), .Y(divider_absoluteValue_B_flipSign_result_20_bF_buf3) );
	BUFX4 BUFX4_666 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_), .Y(divider_absoluteValue_B_flipSign_result_20_bF_buf2) );
	BUFX4 BUFX4_667 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_), .Y(divider_absoluteValue_B_flipSign_result_20_bF_buf1) );
	BUFX4 BUFX4_668 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_), .Y(divider_absoluteValue_B_flipSign_result_20_bF_buf0) );
	BUFX4 BUFX4_669 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .Y(_6627__bF_buf3) );
	BUFX4 BUFX4_670 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .Y(_6627__bF_buf2) );
	BUFX4 BUFX4_671 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .Y(_6627__bF_buf1) );
	BUFX4 BUFX4_672 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .Y(_6627__bF_buf0) );
	BUFX4 BUFX4_673 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf7) );
	BUFX4 BUFX4_674 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf6) );
	BUFX4 BUFX4_675 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf5) );
	BUFX4 BUFX4_676 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf4) );
	BUFX4 BUFX4_677 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf3) );
	BUFX4 BUFX4_678 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf2) );
	BUFX4 BUFX4_679 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf1) );
	BUFX4 BUFX4_680 ( .gnd(gnd), .vdd(vdd), .A(_17392_), .Y(_17392__bF_buf0) );
	BUFX4 BUFX4_681 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_), .Y(aOperand_frameOut_10_bF_buf4) );
	BUFX4 BUFX4_682 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_), .Y(aOperand_frameOut_10_bF_buf3) );
	BUFX4 BUFX4_683 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_), .Y(aOperand_frameOut_10_bF_buf2) );
	BUFX4 BUFX4_684 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_), .Y(aOperand_frameOut_10_bF_buf1) );
	BUFX4 BUFX4_685 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_), .Y(aOperand_frameOut_10_bF_buf0) );
	BUFX4 BUFX4_686 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_), .Y(aOperand_frameOut_5_bF_buf4) );
	BUFX4 BUFX4_687 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_), .Y(aOperand_frameOut_5_bF_buf3) );
	BUFX4 BUFX4_688 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_), .Y(aOperand_frameOut_5_bF_buf2) );
	BUFX4 BUFX4_689 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_), .Y(aOperand_frameOut_5_bF_buf1) );
	BUFX4 BUFX4_690 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_), .Y(aOperand_frameOut_5_bF_buf0) );
	BUFX4 BUFX4_691 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_), .Y(reg_dataIn_23_bF_buf4) );
	BUFX4 BUFX4_692 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_), .Y(reg_dataIn_23_bF_buf3) );
	BUFX4 BUFX4_693 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_), .Y(reg_dataIn_23_bF_buf2) );
	BUFX4 BUFX4_694 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_), .Y(reg_dataIn_23_bF_buf1) );
	BUFX4 BUFX4_695 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_), .Y(reg_dataIn_23_bF_buf0) );
	BUFX4 BUFX4_696 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_), .Y(aOperand_frameOut_0_bF_buf4) );
	BUFX4 BUFX4_697 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_), .Y(aOperand_frameOut_0_bF_buf3) );
	BUFX4 BUFX4_698 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_), .Y(aOperand_frameOut_0_bF_buf2) );
	BUFX4 BUFX4_699 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_), .Y(aOperand_frameOut_0_bF_buf1) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_), .Y(aOperand_frameOut_0_bF_buf0) );
	BUFX4 BUFX4_700 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3255__bF_buf5) );
	BUFX4 BUFX4_701 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3255__bF_buf4) );
	BUFX4 BUFX4_702 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3255__bF_buf3) );
	BUFX4 BUFX4_703 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3255__bF_buf2) );
	BUFX4 BUFX4_704 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3255__bF_buf1) );
	BUFX4 BUFX4_705 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .Y(_3255__bF_buf0) );
	BUFX4 BUFX4_706 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_), .Y(divider_divuResult_21_bF_buf4) );
	BUFX4 BUFX4_707 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_), .Y(divider_divuResult_21_bF_buf3) );
	BUFX4 BUFX4_708 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_), .Y(divider_divuResult_21_bF_buf2) );
	BUFX4 BUFX4_709 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_), .Y(divider_divuResult_21_bF_buf1) );
	BUFX4 BUFX4_710 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_), .Y(divider_divuResult_21_bF_buf0) );
	BUFX4 BUFX4_711 ( .gnd(gnd), .vdd(vdd), .A(_8019_), .Y(_8019__bF_buf3) );
	BUFX4 BUFX4_712 ( .gnd(gnd), .vdd(vdd), .A(_8019_), .Y(_8019__bF_buf2) );
	BUFX4 BUFX4_713 ( .gnd(gnd), .vdd(vdd), .A(_8019_), .Y(_8019__bF_buf1) );
	BUFX4 BUFX4_714 ( .gnd(gnd), .vdd(vdd), .A(_8019_), .Y(_8019__bF_buf0) );
	BUFX4 BUFX4_715 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_), .Y(divider_absoluteValue_B_flipSign_result_18_bF_buf4) );
	BUFX4 BUFX4_716 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_), .Y(divider_absoluteValue_B_flipSign_result_18_bF_buf3) );
	BUFX4 BUFX4_717 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_), .Y(divider_absoluteValue_B_flipSign_result_18_bF_buf2) );
	BUFX4 BUFX4_718 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_), .Y(divider_absoluteValue_B_flipSign_result_18_bF_buf1) );
	BUFX4 BUFX4_719 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_), .Y(divider_absoluteValue_B_flipSign_result_18_bF_buf0) );
	BUFX4 BUFX4_720 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_), .Y(adder_bOperand_16_bF_buf3) );
	BUFX4 BUFX4_721 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_), .Y(adder_bOperand_16_bF_buf2) );
	BUFX4 BUFX4_722 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_), .Y(adder_bOperand_16_bF_buf1) );
	BUFX4 BUFX4_723 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_), .Y(adder_bOperand_16_bF_buf0) );
	BUFX4 BUFX4_724 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_), .Y(reg_dataIn_6_bF_buf4) );
	BUFX4 BUFX4_725 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_), .Y(reg_dataIn_6_bF_buf3) );
	BUFX4 BUFX4_726 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_), .Y(reg_dataIn_6_bF_buf2) );
	BUFX4 BUFX4_727 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_), .Y(reg_dataIn_6_bF_buf1) );
	BUFX4 BUFX4_728 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_), .Y(reg_dataIn_6_bF_buf0) );
	BUFX4 BUFX4_729 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf7) );
	BUFX4 BUFX4_730 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf6) );
	BUFX4 BUFX4_731 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf5) );
	BUFX4 BUFX4_732 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf4) );
	BUFX4 BUFX4_733 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf3) );
	BUFX4 BUFX4_734 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf2) );
	BUFX4 BUFX4_735 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf1) );
	BUFX4 BUFX4_736 ( .gnd(gnd), .vdd(vdd), .A(_19152_), .Y(_19152__bF_buf0) );
	BUFX4 BUFX4_737 ( .gnd(gnd), .vdd(vdd), .A(_20607_), .Y(_20607__bF_buf4) );
	BUFX4 BUFX4_738 ( .gnd(gnd), .vdd(vdd), .A(_20607_), .Y(_20607__bF_buf3) );
	BUFX4 BUFX4_739 ( .gnd(gnd), .vdd(vdd), .A(_20607_), .Y(_20607__bF_buf2) );
	BUFX4 BUFX4_740 ( .gnd(gnd), .vdd(vdd), .A(_20607_), .Y(_20607__bF_buf1) );
	BUFX4 BUFX4_741 ( .gnd(gnd), .vdd(vdd), .A(_20607_), .Y(_20607__bF_buf0) );
	BUFX4 BUFX4_742 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_77__bF_buf4) );
	BUFX4 BUFX4_743 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_77__bF_buf3) );
	BUFX4 BUFX4_744 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_77__bF_buf2) );
	BUFX4 BUFX4_745 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_77__bF_buf1) );
	BUFX4 BUFX4_746 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_77__bF_buf0) );
	BUFX4 BUFX4_747 ( .gnd(gnd), .vdd(vdd), .A(_20595_), .Y(_20595__bF_buf4) );
	BUFX4 BUFX4_748 ( .gnd(gnd), .vdd(vdd), .A(_20595_), .Y(_20595__bF_buf3) );
	BUFX4 BUFX4_749 ( .gnd(gnd), .vdd(vdd), .A(_20595_), .Y(_20595__bF_buf2) );
	BUFX4 BUFX4_750 ( .gnd(gnd), .vdd(vdd), .A(_20595_), .Y(_20595__bF_buf1) );
	BUFX4 BUFX4_751 ( .gnd(gnd), .vdd(vdd), .A(_20595_), .Y(_20595__bF_buf0) );
	BUFX4 BUFX4_752 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_), .Y(divider_absoluteValue_B_flipSign_result_13_bF_buf5) );
	BUFX4 BUFX4_753 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_), .Y(divider_absoluteValue_B_flipSign_result_13_bF_buf4) );
	BUFX4 BUFX4_754 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_), .Y(divider_absoluteValue_B_flipSign_result_13_bF_buf3) );
	BUFX4 BUFX4_755 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_), .Y(divider_absoluteValue_B_flipSign_result_13_bF_buf2) );
	BUFX4 BUFX4_756 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_), .Y(divider_absoluteValue_B_flipSign_result_13_bF_buf1) );
	BUFX4 BUFX4_757 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_), .Y(divider_absoluteValue_B_flipSign_result_13_bF_buf0) );
	BUFX4 BUFX4_758 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .Y(_1983__bF_buf4) );
	BUFX4 BUFX4_759 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .Y(_1983__bF_buf3) );
	BUFX4 BUFX4_760 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .Y(_1983__bF_buf2) );
	BUFX4 BUFX4_761 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .Y(_1983__bF_buf1) );
	BUFX4 BUFX4_762 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .Y(_1983__bF_buf0) );
	BUFX4 BUFX4_763 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2620__bF_buf4) );
	BUFX4 BUFX4_764 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2620__bF_buf3) );
	BUFX4 BUFX4_765 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2620__bF_buf2) );
	BUFX4 BUFX4_766 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2620__bF_buf1) );
	BUFX4 BUFX4_767 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2620__bF_buf0) );
	BUFX4 BUFX4_768 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_), .Y(adder_bOperand_11_bF_buf3) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_), .Y(adder_bOperand_11_bF_buf2) );
	BUFX4 BUFX4_769 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_), .Y(adder_bOperand_11_bF_buf1) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_), .Y(adder_bOperand_11_bF_buf0) );
	BUFX4 BUFX4_770 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_), .Y(reg_dataIn_1_bF_buf4) );
	BUFX4 BUFX4_771 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_), .Y(reg_dataIn_1_bF_buf3) );
	BUFX4 BUFX4_772 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_), .Y(reg_dataIn_1_bF_buf2) );
	BUFX4 BUFX4_773 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_), .Y(reg_dataIn_1_bF_buf1) );
	BUFX4 BUFX4_774 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_), .Y(reg_dataIn_1_bF_buf0) );
	BUFX4 BUFX4_775 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_), .Y(reg_dataIn_16_bF_buf4) );
	BUFX4 BUFX4_776 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_), .Y(reg_dataIn_16_bF_buf3) );
	BUFX4 BUFX4_777 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_), .Y(reg_dataIn_16_bF_buf2) );
	BUFX4 BUFX4_778 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_), .Y(reg_dataIn_16_bF_buf1) );
	BUFX4 BUFX4_779 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_), .Y(reg_dataIn_16_bF_buf0) );
	BUFX4 BUFX4_780 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf7) );
	BUFX4 BUFX4_781 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf6) );
	BUFX4 BUFX4_782 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf5) );
	BUFX4 BUFX4_783 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf4) );
	BUFX4 BUFX4_784 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf3) );
	BUFX4 BUFX4_785 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf2) );
	BUFX4 BUFX4_786 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf1) );
	BUFX4 BUFX4_787 ( .gnd(gnd), .vdd(vdd), .A(_20361_), .Y(_20361__bF_buf0) );
	BUFX4 BUFX4_788 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_), .Y(divider_divuResult_19_bF_buf5) );
	BUFX4 BUFX4_789 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_), .Y(divider_divuResult_19_bF_buf4) );
	BUFX4 BUFX4_790 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_), .Y(divider_divuResult_19_bF_buf3) );
	BUFX4 BUFX4_791 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_), .Y(divider_divuResult_19_bF_buf2) );
	BUFX4 BUFX4_792 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_), .Y(divider_divuResult_19_bF_buf1) );
	BUFX4 BUFX4_793 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_), .Y(divider_divuResult_19_bF_buf0) );
	BUFX4 BUFX4_794 ( .gnd(gnd), .vdd(vdd), .A(_20632_), .Y(_20632__bF_buf4) );
	BUFX4 BUFX4_795 ( .gnd(gnd), .vdd(vdd), .A(_20632_), .Y(_20632__bF_buf3) );
	BUFX4 BUFX4_796 ( .gnd(gnd), .vdd(vdd), .A(_20632_), .Y(_20632__bF_buf2) );
	BUFX4 BUFX4_797 ( .gnd(gnd), .vdd(vdd), .A(_20632_), .Y(_20632__bF_buf1) );
	BUFX4 BUFX4_798 ( .gnd(gnd), .vdd(vdd), .A(_20632_), .Y(_20632__bF_buf0) );
	BUFX4 BUFX4_799 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf6) );
	BUFX4 BUFX4_800 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf5) );
	BUFX4 BUFX4_801 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf4) );
	BUFX4 BUFX4_802 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf3) );
	BUFX4 BUFX4_803 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf2) );
	BUFX4 BUFX4_804 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf1) );
	BUFX4 BUFX4_805 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_), .Y(divider_absoluteValue_B_flipSign_result_6_bF_buf0) );
	BUFX4 BUFX4_806 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf7) );
	BUFX4 BUFX4_807 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf6) );
	BUFX4 BUFX4_808 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf5) );
	BUFX4 BUFX4_809 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf4) );
	BUFX4 BUFX4_810 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf3) );
	BUFX4 BUFX4_811 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf2) );
	BUFX4 BUFX4_812 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf1) );
	BUFX4 BUFX4_813 ( .gnd(gnd), .vdd(vdd), .A(_20590_), .Y(_20590__bF_buf0) );
	BUFX4 BUFX4_814 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_), .Y(adder_bOperand_7_bF_buf5) );
	BUFX4 BUFX4_815 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_), .Y(adder_bOperand_7_bF_buf4) );
	BUFX4 BUFX4_816 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_), .Y(adder_bOperand_7_bF_buf3) );
	BUFX4 BUFX4_817 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_), .Y(adder_bOperand_7_bF_buf2) );
	BUFX4 BUFX4_818 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_), .Y(adder_bOperand_7_bF_buf1) );
	BUFX4 BUFX4_819 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_), .Y(adder_bOperand_7_bF_buf0) );
	BUFX4 BUFX4_820 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_), .Y(reg_dataIn_11_bF_buf4) );
	BUFX4 BUFX4_821 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_), .Y(reg_dataIn_11_bF_buf3) );
	BUFX4 BUFX4_822 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_), .Y(reg_dataIn_11_bF_buf2) );
	BUFX4 BUFX4_823 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_), .Y(reg_dataIn_11_bF_buf1) );
	BUFX4 BUFX4_824 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_), .Y(reg_dataIn_11_bF_buf0) );
	BUFX4 BUFX4_825 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_), .Y(divider_divuResult_14_bF_buf4) );
	BUFX4 BUFX4_826 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_), .Y(divider_divuResult_14_bF_buf3) );
	BUFX4 BUFX4_827 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_), .Y(divider_divuResult_14_bF_buf2) );
	BUFX4 BUFX4_828 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_), .Y(divider_divuResult_14_bF_buf1) );
	BUFX4 BUFX4_829 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_), .Y(divider_divuResult_14_bF_buf0) );
	BUFX4 BUFX4_830 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf7) );
	BUFX4 BUFX4_831 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf6) );
	BUFX4 BUFX4_832 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf5) );
	BUFX4 BUFX4_833 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf4) );
	BUFX4 BUFX4_834 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf3) );
	BUFX4 BUFX4_835 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf2) );
	BUFX4 BUFX4_836 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf1) );
	BUFX4 BUFX4_837 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_), .Y(divider_absoluteValue_B_flipSign_result_1_bF_buf0) );
	BUFX4 BUFX4_838 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_), .Y(adder_bOperand_2_bF_buf5) );
	BUFX4 BUFX4_839 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_), .Y(adder_bOperand_2_bF_buf4) );
	BUFX4 BUFX4_840 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_), .Y(adder_bOperand_2_bF_buf3) );
	BUFX4 BUFX4_841 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_), .Y(adder_bOperand_2_bF_buf2) );
	BUFX4 BUFX4_842 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_), .Y(adder_bOperand_2_bF_buf1) );
	BUFX4 BUFX4_843 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_), .Y(adder_bOperand_2_bF_buf0) );
	BUFX4 BUFX4_844 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_435__bF_buf5) );
	BUFX4 BUFX4_845 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_435__bF_buf4) );
	BUFX4 BUFX4_846 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_435__bF_buf3) );
	BUFX4 BUFX4_847 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_435__bF_buf2) );
	BUFX4 BUFX4_848 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_435__bF_buf1) );
	BUFX4 BUFX4_849 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_435__bF_buf0) );
	BUFX4 BUFX4_850 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .Y(_3171__bF_buf3) );
	BUFX4 BUFX4_851 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .Y(_3171__bF_buf2) );
	BUFX4 BUFX4_852 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .Y(_3171__bF_buf1) );
	BUFX4 BUFX4_853 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .Y(_3171__bF_buf0) );
	BUFX4 BUFX4_854 ( .gnd(gnd), .vdd(vdd), .A(_20588_), .Y(_20588__bF_buf5) );
	BUFX4 BUFX4_855 ( .gnd(gnd), .vdd(vdd), .A(_20588_), .Y(_20588__bF_buf4) );
	BUFX4 BUFX4_856 ( .gnd(gnd), .vdd(vdd), .A(_20588_), .Y(_20588__bF_buf3) );
	BUFX4 BUFX4_857 ( .gnd(gnd), .vdd(vdd), .A(_20588_), .Y(_20588__bF_buf2) );
	BUFX4 BUFX4_858 ( .gnd(gnd), .vdd(vdd), .A(_20588_), .Y(_20588__bF_buf1) );
	BUFX4 BUFX4_859 ( .gnd(gnd), .vdd(vdd), .A(_20588_), .Y(_20588__bF_buf0) );
	BUFX4 BUFX4_860 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf6) );
	BUFX4 BUFX4_861 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf5) );
	BUFX4 BUFX4_862 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf4) );
	BUFX4 BUFX4_863 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf3) );
	BUFX4 BUFX4_864 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf2) );
	BUFX4 BUFX4_865 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf1) );
	BUFX4 BUFX4_866 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_), .Y(divider_divuResult_5_bF_buf0) );
	BUFX4 BUFX4_867 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .Y(_1615__bF_buf4) );
	BUFX4 BUFX4_868 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .Y(_1615__bF_buf3) );
	BUFX4 BUFX4_869 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .Y(_1615__bF_buf2) );
	BUFX4 BUFX4_870 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .Y(_1615__bF_buf1) );
	BUFX4 BUFX4_871 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .Y(_1615__bF_buf0) );
	BUFX4 BUFX4_872 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2240__bF_buf4) );
	BUFX4 BUFX4_873 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2240__bF_buf3) );
	BUFX4 BUFX4_874 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2240__bF_buf2) );
	BUFX4 BUFX4_875 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2240__bF_buf1) );
	BUFX4 BUFX4_876 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2240__bF_buf0) );
	BUFX4 BUFX4_877 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf6) );
	BUFX4 BUFX4_878 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf5) );
	BUFX4 BUFX4_879 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf4) );
	BUFX4 BUFX4_880 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf3) );
	BUFX4 BUFX4_881 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf2) );
	BUFX4 BUFX4_882 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf1) );
	BUFX4 BUFX4_883 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .Y(_8664__bF_buf0) );
	BUFX4 BUFX4_884 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf3) );
	BUFX4 BUFX4_885 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf2) );
	BUFX4 BUFX4_886 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf1) );
	BUFX4 BUFX4_887 ( .gnd(gnd), .vdd(vdd), .A(_8062_), .Y(_8062__bF_buf0) );
	BUFX4 BUFX4_888 ( .gnd(gnd), .vdd(vdd), .A(_17373_), .Y(_17373__bF_buf5) );
	BUFX4 BUFX4_889 ( .gnd(gnd), .vdd(vdd), .A(_17373_), .Y(_17373__bF_buf4) );
	BUFX4 BUFX4_890 ( .gnd(gnd), .vdd(vdd), .A(_17373_), .Y(_17373__bF_buf3) );
	BUFX4 BUFX4_891 ( .gnd(gnd), .vdd(vdd), .A(_17373_), .Y(_17373__bF_buf2) );
	BUFX4 BUFX4_892 ( .gnd(gnd), .vdd(vdd), .A(_17373_), .Y(_17373__bF_buf1) );
	BUFX4 BUFX4_893 ( .gnd(gnd), .vdd(vdd), .A(_17373_), .Y(_17373__bF_buf0) );
	BUFX4 BUFX4_894 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf6) );
	BUFX4 BUFX4_895 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf5) );
	BUFX4 BUFX4_896 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf4) );
	BUFX4 BUFX4_897 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf3) );
	BUFX4 BUFX4_898 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf2) );
	BUFX4 BUFX4_899 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf1) );
	BUFX4 BUFX4_900 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_), .Y(divider_divuResult_0_bF_buf0) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_), .Y(aOperand_frameOut_21_bF_buf4) );
	BUFX4 BUFX4_901 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_), .Y(aOperand_frameOut_21_bF_buf3) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_), .Y(aOperand_frameOut_21_bF_buf2) );
	BUFX4 BUFX4_902 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_), .Y(aOperand_frameOut_21_bF_buf1) );
	BUFX4 BUFX4_903 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_), .Y(aOperand_frameOut_21_bF_buf0) );
	BUFX4 BUFX4_904 ( .gnd(gnd), .vdd(vdd), .A(_17440_), .Y(_17440__bF_buf4) );
	BUFX4 BUFX4_905 ( .gnd(gnd), .vdd(vdd), .A(_17440_), .Y(_17440__bF_buf3) );
	BUFX4 BUFX4_906 ( .gnd(gnd), .vdd(vdd), .A(_17440_), .Y(_17440__bF_buf2) );
	BUFX4 BUFX4_907 ( .gnd(gnd), .vdd(vdd), .A(_17440_), .Y(_17440__bF_buf1) );
	BUFX4 BUFX4_908 ( .gnd(gnd), .vdd(vdd), .A(_17440_), .Y(_17440__bF_buf0) );
	BUFX4 BUFX4_909 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .Y(_4065__bF_buf4) );
	BUFX4 BUFX4_910 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .Y(_4065__bF_buf3) );
	BUFX4 BUFX4_911 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .Y(_4065__bF_buf2) );
	BUFX4 BUFX4_912 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .Y(_4065__bF_buf1) );
	BUFX4 BUFX4_913 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .Y(_4065__bF_buf0) );
	BUFX4 BUFX4_914 ( .gnd(gnd), .vdd(vdd), .A(_15812_), .Y(_15812__bF_buf3) );
	BUFX4 BUFX4_915 ( .gnd(gnd), .vdd(vdd), .A(_15812_), .Y(_15812__bF_buf2) );
	BUFX4 BUFX4_916 ( .gnd(gnd), .vdd(vdd), .A(_15812_), .Y(_15812__bF_buf1) );
	BUFX4 BUFX4_917 ( .gnd(gnd), .vdd(vdd), .A(_15812_), .Y(_15812__bF_buf0) );
	BUFX4 BUFX4_918 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf7) );
	BUFX4 BUFX4_919 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf6) );
	BUFX4 BUFX4_920 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf5) );
	BUFX4 BUFX4_921 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf4) );
	BUFX4 BUFX4_922 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf3) );
	BUFX4 BUFX4_923 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf2) );
	BUFX4 BUFX4_924 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf1) );
	BUFX4 BUFX4_925 ( .gnd(gnd), .vdd(vdd), .A(_19499_), .Y(_19499__bF_buf0) );
	BUFX4 BUFX4_926 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf7) );
	BUFX4 BUFX4_927 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf6) );
	BUFX4 BUFX4_928 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf5) );
	BUFX4 BUFX4_929 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf4) );
	BUFX4 BUFX4_930 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf3) );
	BUFX4 BUFX4_931 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf2) );
	BUFX4 BUFX4_932 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf1) );
	BUFX4 BUFX4_933 ( .gnd(gnd), .vdd(vdd), .A(_19668_), .Y(_19668__bF_buf0) );
	BUFX4 BUFX4_934 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_), .Y(aOperand_frameOut_19_bF_buf4) );
	BUFX4 BUFX4_935 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_), .Y(aOperand_frameOut_19_bF_buf3) );
	BUFX4 BUFX4_936 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_), .Y(aOperand_frameOut_19_bF_buf2) );
	BUFX4 BUFX4_937 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_), .Y(aOperand_frameOut_19_bF_buf1) );
	BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_), .Y(aOperand_frameOut_19_bF_buf0) );
	BUFX4 BUFX4_938 ( .gnd(gnd), .vdd(vdd), .A(_3261_), .Y(_3261__bF_buf3) );
	BUFX4 BUFX4_939 ( .gnd(gnd), .vdd(vdd), .A(_3261_), .Y(_3261__bF_buf2) );
	BUFX4 BUFX4_940 ( .gnd(gnd), .vdd(vdd), .A(_3261_), .Y(_3261__bF_buf1) );
	BUFX4 BUFX4_941 ( .gnd(gnd), .vdd(vdd), .A(_3261_), .Y(_3261__bF_buf0) );
	BUFX4 BUFX4_942 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf7) );
	BUFX4 BUFX4_943 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf6) );
	BUFX4 BUFX4_944 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf5) );
	BUFX4 BUFX4_945 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf4) );
	BUFX4 BUFX4_946 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf3) );
	BUFX4 BUFX4_947 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf2) );
	BUFX4 BUFX4_948 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf1) );
	BUFX4 BUFX4_949 ( .gnd(gnd), .vdd(vdd), .A(_19837_), .Y(_19837__bF_buf0) );
	BUFX4 BUFX4_950 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .Y(_10678__bF_buf5) );
	BUFX4 BUFX4_951 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .Y(_10678__bF_buf4) );
	BUFX4 BUFX4_952 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .Y(_10678__bF_buf3) );
	BUFX4 BUFX4_953 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .Y(_10678__bF_buf2) );
	BUFX4 BUFX4_954 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .Y(_10678__bF_buf1) );
	BUFX4 BUFX4_955 ( .gnd(gnd), .vdd(vdd), .A(_10678_), .Y(_10678__bF_buf0) );
	BUFX4 BUFX4_956 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .Y(_1265__bF_buf5) );
	BUFX4 BUFX4_957 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .Y(_1265__bF_buf4) );
	BUFX4 BUFX4_958 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .Y(_1265__bF_buf3) );
	BUFX4 BUFX4_959 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .Y(_1265__bF_buf2) );
	BUFX4 BUFX4_960 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .Y(_1265__bF_buf1) );
	BUFX4 BUFX4_961 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .Y(_1265__bF_buf0) );
	BUFX4 BUFX4_962 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .Y(_1494__bF_buf4) );
	BUFX4 BUFX4_963 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .Y(_1494__bF_buf3) );
	BUFX4 BUFX4_964 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .Y(_1494__bF_buf2) );
	BUFX4 BUFX4_965 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .Y(_1494__bF_buf1) );
	BUFX4 BUFX4_966 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .Y(_1494__bF_buf0) );
	BUFX4 BUFX4_967 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf7) );
	BUFX4 BUFX4_968 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf6) );
	BUFX4 BUFX4_969 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf5) );
	BUFX4 BUFX4_970 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf4) );
	BUFX4 BUFX4_971 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf3) );
	BUFX4 BUFX4_972 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf2) );
	BUFX4 BUFX4_973 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf1) );
	BUFX4 BUFX4_974 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut), .Y(immediateSelect_frameOut_bF_buf0) );
	BUFX4 BUFX4_975 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf7) );
	BUFX4 BUFX4_976 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf6) );
	BUFX4 BUFX4_977 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf5) );
	BUFX4 BUFX4_978 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf4) );
	BUFX4 BUFX4_979 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf3) );
	BUFX4 BUFX4_980 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf2) );
	BUFX4 BUFX4_981 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf1) );
	BUFX4 BUFX4_982 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf0) );
	BUFX4 BUFX4_983 ( .gnd(gnd), .vdd(vdd), .A(_17408_), .Y(_17408__bF_buf4) );
	BUFX4 BUFX4_984 ( .gnd(gnd), .vdd(vdd), .A(_17408_), .Y(_17408__bF_buf3) );
	BUFX4 BUFX4_985 ( .gnd(gnd), .vdd(vdd), .A(_17408_), .Y(_17408__bF_buf2) );
	BUFX4 BUFX4_986 ( .gnd(gnd), .vdd(vdd), .A(_17408_), .Y(_17408__bF_buf1) );
	BUFX4 BUFX4_987 ( .gnd(gnd), .vdd(vdd), .A(_17408_), .Y(_17408__bF_buf0) );
	BUFX4 BUFX4_988 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_), .Y(divider_absoluteValue_B_flipSign_result_24_bF_buf3) );
	BUFX4 BUFX4_989 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_), .Y(divider_absoluteValue_B_flipSign_result_24_bF_buf2) );
	BUFX4 BUFX4_990 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_), .Y(divider_absoluteValue_B_flipSign_result_24_bF_buf1) );
	BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_), .Y(divider_absoluteValue_B_flipSign_result_24_bF_buf0) );
	BUFX4 BUFX4_991 ( .gnd(gnd), .vdd(vdd), .A(_20576_), .Y(_20576__bF_buf4) );
	BUFX4 BUFX4_992 ( .gnd(gnd), .vdd(vdd), .A(_20576_), .Y(_20576__bF_buf3) );
	BUFX4 BUFX4_993 ( .gnd(gnd), .vdd(vdd), .A(_20576_), .Y(_20576__bF_buf2) );
	BUFX4 BUFX4_994 ( .gnd(gnd), .vdd(vdd), .A(_20576_), .Y(_20576__bF_buf1) );
	BUFX4 BUFX4_995 ( .gnd(gnd), .vdd(vdd), .A(_20576_), .Y(_20576__bF_buf0) );
	BUFX4 BUFX4_996 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf7) );
	BUFX4 BUFX4_997 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf6) );
	BUFX4 BUFX4_998 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf5) );
	BUFX4 BUFX4_999 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf4) );
	BUFX4 BUFX4_1000 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf3) );
	BUFX4 BUFX4_1001 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf2) );
	BUFX4 BUFX4_1002 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf1) );
	BUFX4 BUFX4_1003 ( .gnd(gnd), .vdd(vdd), .A(_19362_), .Y(_19362__bF_buf0) );
	BUFX4 BUFX4_1004 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf7) );
	BUFX4 BUFX4_1005 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf6) );
	BUFX4 BUFX4_1006 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf5) );
	BUFX4 BUFX4_1007 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf4) );
	BUFX4 BUFX4_1008 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf3) );
	BUFX4 BUFX4_1009 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf2) );
	BUFX4 BUFX4_1010 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf1) );
	BUFX4 BUFX4_1011 ( .gnd(gnd), .vdd(vdd), .A(_19904_), .Y(_19904__bF_buf0) );
	BUFX4 BUFX4_1012 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_), .Y(adder_bOperand_22_bF_buf3) );
	BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_), .Y(adder_bOperand_22_bF_buf2) );
	BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_), .Y(adder_bOperand_22_bF_buf1) );
	BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_), .Y(adder_bOperand_22_bF_buf0) );
	BUFX4 BUFX4_1013 ( .gnd(gnd), .vdd(vdd), .A(_17306_), .Y(_17306__bF_buf3) );
	BUFX4 BUFX4_1014 ( .gnd(gnd), .vdd(vdd), .A(_17306_), .Y(_17306__bF_buf2) );
	BUFX4 BUFX4_1015 ( .gnd(gnd), .vdd(vdd), .A(_17306_), .Y(_17306__bF_buf1) );
	BUFX4 BUFX4_1016 ( .gnd(gnd), .vdd(vdd), .A(_17306_), .Y(_17306__bF_buf0) );
	BUFX4 BUFX4_1017 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_), .Y(aOperand_frameOut_14_bF_buf4) );
	BUFX4 BUFX4_1018 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_), .Y(aOperand_frameOut_14_bF_buf3) );
	BUFX4 BUFX4_1019 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_), .Y(aOperand_frameOut_14_bF_buf2) );
	BUFX4 BUFX4_1020 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_), .Y(aOperand_frameOut_14_bF_buf1) );
	BUFX4 BUFX4_1021 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_), .Y(aOperand_frameOut_14_bF_buf0) );
	BUFX4 BUFX4_1022 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_), .Y(aOperand_frameOut_9_bF_buf4) );
	BUFX4 BUFX4_1023 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_), .Y(aOperand_frameOut_9_bF_buf3) );
	BUFX4 BUFX4_1024 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_), .Y(aOperand_frameOut_9_bF_buf2) );
	BUFX4 BUFX4_1025 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_), .Y(aOperand_frameOut_9_bF_buf1) );
	BUFX4 BUFX4_1026 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_), .Y(aOperand_frameOut_9_bF_buf0) );
	BUFX4 BUFX4_1027 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_), .Y(reg_dataIn_27_bF_buf4) );
	BUFX4 BUFX4_1028 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_), .Y(reg_dataIn_27_bF_buf3) );
	BUFX4 BUFX4_1029 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_), .Y(reg_dataIn_27_bF_buf2) );
	BUFX4 BUFX4_1030 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_), .Y(reg_dataIn_27_bF_buf1) );
	BUFX4 BUFX4_1031 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_), .Y(reg_dataIn_27_bF_buf0) );
	BUFX4 BUFX4_1032 ( .gnd(gnd), .vdd(vdd), .A(_17433_), .Y(_17433__bF_buf4) );
	BUFX4 BUFX4_1033 ( .gnd(gnd), .vdd(vdd), .A(_17433_), .Y(_17433__bF_buf3) );
	BUFX4 BUFX4_1034 ( .gnd(gnd), .vdd(vdd), .A(_17433_), .Y(_17433__bF_buf2) );
	BUFX4 BUFX4_1035 ( .gnd(gnd), .vdd(vdd), .A(_17433_), .Y(_17433__bF_buf1) );
	BUFX4 BUFX4_1036 ( .gnd(gnd), .vdd(vdd), .A(_17433_), .Y(_17433__bF_buf0) );
	BUFX4 BUFX4_1037 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_83__bF_buf4) );
	BUFX4 BUFX4_1038 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_83__bF_buf3) );
	BUFX4 BUFX4_1039 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_83__bF_buf2) );
	BUFX4 BUFX4_1040 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_83__bF_buf1) );
	BUFX4 BUFX4_1041 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_83__bF_buf0) );
	BUFX4 BUFX4_1042 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_), .Y(aOperand_frameOut_4_bF_buf4) );
	BUFX4 BUFX4_1043 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_), .Y(aOperand_frameOut_4_bF_buf3) );
	BUFX4 BUFX4_1044 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_), .Y(aOperand_frameOut_4_bF_buf2) );
	BUFX4 BUFX4_1045 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_), .Y(aOperand_frameOut_4_bF_buf1) );
	BUFX4 BUFX4_1046 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_), .Y(aOperand_frameOut_4_bF_buf0) );
	BUFX4 BUFX4_1047 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_), .Y(reg_dataIn_22_bF_buf4) );
	BUFX4 BUFX4_1048 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_), .Y(reg_dataIn_22_bF_buf3) );
	BUFX4 BUFX4_1049 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_), .Y(reg_dataIn_22_bF_buf2) );
	BUFX4 BUFX4_1050 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_), .Y(reg_dataIn_22_bF_buf1) );
	BUFX4 BUFX4_1051 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_), .Y(reg_dataIn_22_bF_buf0) );
	BUFX4 BUFX4_1052 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .Y(_7450__bF_buf5) );
	BUFX4 BUFX4_1053 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .Y(_7450__bF_buf4) );
	BUFX4 BUFX4_1054 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .Y(_7450__bF_buf3) );
	BUFX4 BUFX4_1055 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .Y(_7450__bF_buf2) );
	BUFX4 BUFX4_1056 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .Y(_7450__bF_buf1) );
	BUFX4 BUFX4_1057 ( .gnd(gnd), .vdd(vdd), .A(_7450_), .Y(_7450__bF_buf0) );
	BUFX4 BUFX4_1058 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .Y(_3789__bF_buf4) );
	BUFX4 BUFX4_1059 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .Y(_3789__bF_buf3) );
	BUFX4 BUFX4_1060 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .Y(_3789__bF_buf2) );
	BUFX4 BUFX4_1061 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .Y(_3789__bF_buf1) );
	BUFX4 BUFX4_1062 ( .gnd(gnd), .vdd(vdd), .A(_3789_), .Y(_3789__bF_buf0) );
	BUFX4 BUFX4_1063 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .Y(_13436__bF_buf3) );
	BUFX4 BUFX4_1064 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .Y(_13436__bF_buf2) );
	BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .Y(_13436__bF_buf1) );
	BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_13436_), .Y(_13436__bF_buf0) );
	BUFX4 BUFX4_1065 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_), .Y(divider_divuResult_20_bF_buf3) );
	BUFX4 BUFX4_1066 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_), .Y(divider_divuResult_20_bF_buf2) );
	BUFX4 BUFX4_1067 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_), .Y(divider_divuResult_20_bF_buf1) );
	BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_), .Y(divider_divuResult_20_bF_buf0) );
	BUFX4 BUFX4_1068 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_), .Y(divider_absoluteValue_B_flipSign_result_17_bF_buf4) );
	BUFX4 BUFX4_1069 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_), .Y(divider_absoluteValue_B_flipSign_result_17_bF_buf3) );
	BUFX4 BUFX4_1070 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_), .Y(divider_absoluteValue_B_flipSign_result_17_bF_buf2) );
	BUFX4 BUFX4_1071 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_), .Y(divider_absoluteValue_B_flipSign_result_17_bF_buf1) );
	BUFX4 BUFX4_1072 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_), .Y(divider_absoluteValue_B_flipSign_result_17_bF_buf0) );
	BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_), .Y(adder_bOperand_15_bF_buf4) );
	BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_), .Y(adder_bOperand_15_bF_buf3) );
	BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_), .Y(adder_bOperand_15_bF_buf2) );
	BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_), .Y(adder_bOperand_15_bF_buf1) );
	BUFX4 BUFX4_1073 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_), .Y(adder_bOperand_15_bF_buf0) );
	BUFX4 BUFX4_1074 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf7) );
	BUFX4 BUFX4_1075 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf6) );
	BUFX4 BUFX4_1076 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf5) );
	BUFX4 BUFX4_1077 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf4) );
	BUFX4 BUFX4_1078 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf3) );
	BUFX4 BUFX4_1079 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf2) );
	BUFX4 BUFX4_1080 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf1) );
	BUFX4 BUFX4_1081 ( .gnd(gnd), .vdd(vdd), .A(_20166_), .Y(_20166__bF_buf0) );
	BUFX4 BUFX4_1082 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_), .Y(reg_dataIn_5_bF_buf4) );
	BUFX4 BUFX4_1083 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_), .Y(reg_dataIn_5_bF_buf3) );
	BUFX4 BUFX4_1084 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_), .Y(reg_dataIn_5_bF_buf2) );
	BUFX4 BUFX4_1085 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_), .Y(reg_dataIn_5_bF_buf1) );
	BUFX4 BUFX4_1086 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_), .Y(reg_dataIn_5_bF_buf0) );
	BUFX4 BUFX4_1087 ( .gnd(gnd), .vdd(vdd), .A(_20606_), .Y(_20606__bF_buf4) );
	BUFX4 BUFX4_1088 ( .gnd(gnd), .vdd(vdd), .A(_20606_), .Y(_20606__bF_buf3) );
	BUFX4 BUFX4_1089 ( .gnd(gnd), .vdd(vdd), .A(_20606_), .Y(_20606__bF_buf2) );
	BUFX4 BUFX4_1090 ( .gnd(gnd), .vdd(vdd), .A(_20606_), .Y(_20606__bF_buf1) );
	BUFX4 BUFX4_1091 ( .gnd(gnd), .vdd(vdd), .A(_20606_), .Y(_20606__bF_buf0) );
	BUFX4 BUFX4_1092 ( .gnd(gnd), .vdd(vdd), .A(_17456_), .Y(_17456__bF_buf4) );
	BUFX4 BUFX4_1093 ( .gnd(gnd), .vdd(vdd), .A(_17456_), .Y(_17456__bF_buf3) );
	BUFX4 BUFX4_1094 ( .gnd(gnd), .vdd(vdd), .A(_17456_), .Y(_17456__bF_buf2) );
	BUFX4 BUFX4_1095 ( .gnd(gnd), .vdd(vdd), .A(_17456_), .Y(_17456__bF_buf1) );
	BUFX4 BUFX4_1096 ( .gnd(gnd), .vdd(vdd), .A(_17456_), .Y(_17456__bF_buf0) );
	BUFX4 BUFX4_1097 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf6) );
	BUFX4 BUFX4_1098 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf5) );
	BUFX4 BUFX4_1099 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf4) );
	BUFX4 BUFX4_1100 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf3) );
	BUFX4 BUFX4_1101 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf2) );
	BUFX4 BUFX4_1102 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf1) );
	BUFX4 BUFX4_1103 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_), .Y(aLoc_frameOut_4_bF_buf0) );
	BUFX4 BUFX4_1104 ( .gnd(gnd), .vdd(vdd), .A(_20594_), .Y(_20594__bF_buf4) );
	BUFX4 BUFX4_1105 ( .gnd(gnd), .vdd(vdd), .A(_20594_), .Y(_20594__bF_buf3) );
	BUFX4 BUFX4_1106 ( .gnd(gnd), .vdd(vdd), .A(_20594_), .Y(_20594__bF_buf2) );
	BUFX4 BUFX4_1107 ( .gnd(gnd), .vdd(vdd), .A(_20594_), .Y(_20594__bF_buf1) );
	BUFX4 BUFX4_1108 ( .gnd(gnd), .vdd(vdd), .A(_20594_), .Y(_20594__bF_buf0) );
	BUFX4 BUFX4_1109 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_), .Y(divider_absoluteValue_B_flipSign_result_12_bF_buf5) );
	BUFX4 BUFX4_1110 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_), .Y(divider_absoluteValue_B_flipSign_result_12_bF_buf4) );
	BUFX4 BUFX4_1111 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_), .Y(divider_absoluteValue_B_flipSign_result_12_bF_buf3) );
	BUFX4 BUFX4_1112 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_), .Y(divider_absoluteValue_B_flipSign_result_12_bF_buf2) );
	BUFX4 BUFX4_1113 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_), .Y(divider_absoluteValue_B_flipSign_result_12_bF_buf1) );
	BUFX4 BUFX4_1114 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_), .Y(divider_absoluteValue_B_flipSign_result_12_bF_buf0) );
	BUFX4 BUFX4_1115 ( .gnd(gnd), .vdd(vdd), .A(_17384_), .Y(_17384__bF_buf4) );
	BUFX4 BUFX4_1116 ( .gnd(gnd), .vdd(vdd), .A(_17384_), .Y(_17384__bF_buf3) );
	BUFX4 BUFX4_1117 ( .gnd(gnd), .vdd(vdd), .A(_17384_), .Y(_17384__bF_buf2) );
	BUFX4 BUFX4_1118 ( .gnd(gnd), .vdd(vdd), .A(_17384_), .Y(_17384__bF_buf1) );
	BUFX4 BUFX4_1119 ( .gnd(gnd), .vdd(vdd), .A(_17384_), .Y(_17384__bF_buf0) );
	BUFX4 BUFX4_1120 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_), .Y(adder_bOperand_10_bF_buf4) );
	BUFX4 BUFX4_1121 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_), .Y(adder_bOperand_10_bF_buf3) );
	BUFX4 BUFX4_1122 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_), .Y(adder_bOperand_10_bF_buf2) );
	BUFX4 BUFX4_1123 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_), .Y(adder_bOperand_10_bF_buf1) );
	BUFX4 BUFX4_1124 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_), .Y(adder_bOperand_10_bF_buf0) );
	BUFX4 BUFX4_1125 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf7) );
	BUFX4 BUFX4_1126 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf6) );
	BUFX4 BUFX4_1127 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf5) );
	BUFX4 BUFX4_1128 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf4) );
	BUFX4 BUFX4_1129 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf3) );
	BUFX4 BUFX4_1130 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf2) );
	BUFX4 BUFX4_1131 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf1) );
	BUFX4 BUFX4_1132 ( .gnd(gnd), .vdd(vdd), .A(_20492_), .Y(_20492__bF_buf0) );
	BUFX4 BUFX4_1133 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_), .Y(reg_dataIn_0_bF_buf4) );
	BUFX4 BUFX4_1134 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_), .Y(reg_dataIn_0_bF_buf3) );
	BUFX4 BUFX4_1135 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_), .Y(reg_dataIn_0_bF_buf2) );
	BUFX4 BUFX4_1136 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_), .Y(reg_dataIn_0_bF_buf1) );
	BUFX4 BUFX4_1137 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_), .Y(reg_dataIn_0_bF_buf0) );
	BUFX4 BUFX4_1138 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf7) );
	BUFX4 BUFX4_1139 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf6) );
	BUFX4 BUFX4_1140 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf5) );
	BUFX4 BUFX4_1141 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf4) );
	BUFX4 BUFX4_1142 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf3) );
	BUFX4 BUFX4_1143 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf2) );
	BUFX4 BUFX4_1144 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf1) );
	BUFX4 BUFX4_1145 ( .gnd(gnd), .vdd(vdd), .A(_20101_), .Y(_20101__bF_buf0) );
	BUFX4 BUFX4_1146 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_), .Y(reg_dataIn_15_bF_buf4) );
	BUFX4 BUFX4_1147 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_), .Y(reg_dataIn_15_bF_buf3) );
	BUFX4 BUFX4_1148 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_), .Y(reg_dataIn_15_bF_buf2) );
	BUFX4 BUFX4_1149 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_), .Y(reg_dataIn_15_bF_buf1) );
	BUFX4 BUFX4_1150 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_), .Y(reg_dataIn_15_bF_buf0) );
	BUFX4 BUFX4_1151 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_), .Y(divider_divuResult_18_bF_buf5) );
	BUFX4 BUFX4_1152 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_), .Y(divider_divuResult_18_bF_buf4) );
	BUFX4 BUFX4_1153 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_), .Y(divider_divuResult_18_bF_buf3) );
	BUFX4 BUFX4_1154 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_), .Y(divider_divuResult_18_bF_buf2) );
	BUFX4 BUFX4_1155 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_), .Y(divider_divuResult_18_bF_buf1) );
	BUFX4 BUFX4_1156 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_), .Y(divider_divuResult_18_bF_buf0) );
	BUFX4 BUFX4_1157 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf7) );
	BUFX4 BUFX4_1158 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf6) );
	BUFX4 BUFX4_1159 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf5) );
	BUFX4 BUFX4_1160 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf4) );
	BUFX4 BUFX4_1161 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf3) );
	BUFX4 BUFX4_1162 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf2) );
	BUFX4 BUFX4_1163 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf1) );
	BUFX4 BUFX4_1164 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_), .Y(divider_absoluteValue_B_flipSign_result_5_bF_buf0) );
	BUFX4 BUFX4_1165 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf6) );
	BUFX4 BUFX4_1166 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf5) );
	BUFX4 BUFX4_1167 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf4) );
	BUFX4 BUFX4_1168 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf3) );
	BUFX4 BUFX4_1169 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf2) );
	BUFX4 BUFX4_1170 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf1) );
	BUFX4 BUFX4_1171 ( .gnd(gnd), .vdd(vdd), .A(_8971_), .Y(_8971__bF_buf0) );
	BUFX4 BUFX4_1172 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_71__bF_buf4) );
	BUFX4 BUFX4_1173 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_71__bF_buf3) );
	BUFX4 BUFX4_1174 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_71__bF_buf2) );
	BUFX4 BUFX4_1175 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_71__bF_buf1) );
	BUFX4 BUFX4_1176 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_71__bF_buf0) );
	BUFX4 BUFX4_1177 ( .gnd(gnd), .vdd(vdd), .A(_14728_), .Y(_14728__bF_buf3) );
	BUFX4 BUFX4_1178 ( .gnd(gnd), .vdd(vdd), .A(_14728_), .Y(_14728__bF_buf2) );
	BUFX4 BUFX4_1179 ( .gnd(gnd), .vdd(vdd), .A(_14728_), .Y(_14728__bF_buf1) );
	BUFX4 BUFX4_1180 ( .gnd(gnd), .vdd(vdd), .A(_14728_), .Y(_14728__bF_buf0) );
	BUFX4 BUFX4_1181 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_), .Y(adder_bOperand_6_bF_buf5) );
	BUFX4 BUFX4_1182 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_), .Y(adder_bOperand_6_bF_buf4) );
	BUFX4 BUFX4_1183 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_), .Y(adder_bOperand_6_bF_buf3) );
	BUFX4 BUFX4_1184 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_), .Y(adder_bOperand_6_bF_buf2) );
	BUFX4 BUFX4_1185 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_), .Y(adder_bOperand_6_bF_buf1) );
	BUFX4 BUFX4_1186 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_), .Y(adder_bOperand_6_bF_buf0) );
	BUFX4 BUFX4_1187 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_), .Y(reg_dataIn_10_bF_buf4) );
	BUFX4 BUFX4_1188 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_), .Y(reg_dataIn_10_bF_buf3) );
	BUFX4 BUFX4_1189 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_), .Y(reg_dataIn_10_bF_buf2) );
	BUFX4 BUFX4_1190 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_), .Y(reg_dataIn_10_bF_buf1) );
	BUFX4 BUFX4_1191 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_), .Y(reg_dataIn_10_bF_buf0) );
	BUFX4 BUFX4_1192 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_), .Y(divider_divuResult_13_bF_buf5) );
	BUFX4 BUFX4_1193 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_), .Y(divider_divuResult_13_bF_buf4) );
	BUFX4 BUFX4_1194 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_), .Y(divider_divuResult_13_bF_buf3) );
	BUFX4 BUFX4_1195 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_), .Y(divider_divuResult_13_bF_buf2) );
	BUFX4 BUFX4_1196 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_), .Y(divider_divuResult_13_bF_buf1) );
	BUFX4 BUFX4_1197 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_), .Y(divider_divuResult_13_bF_buf0) );
	BUFX4 BUFX4_1198 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_), .Y(divider_absoluteValue_B_flipSign_result_0_bF_buf5) );
	BUFX4 BUFX4_1199 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_), .Y(divider_absoluteValue_B_flipSign_result_0_bF_buf4) );
	BUFX4 BUFX4_1200 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_), .Y(divider_absoluteValue_B_flipSign_result_0_bF_buf3) );
	BUFX4 BUFX4_1201 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_), .Y(divider_absoluteValue_B_flipSign_result_0_bF_buf2) );
	BUFX4 BUFX4_1202 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_), .Y(divider_absoluteValue_B_flipSign_result_0_bF_buf1) );
	BUFX4 BUFX4_1203 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_), .Y(divider_absoluteValue_B_flipSign_result_0_bF_buf0) );
	BUFX4 BUFX4_1204 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf6) );
	BUFX4 BUFX4_1205 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf5) );
	BUFX4 BUFX4_1206 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf4) );
	BUFX4 BUFX4_1207 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf3) );
	BUFX4 BUFX4_1208 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf2) );
	BUFX4 BUFX4_1209 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf1) );
	BUFX4 BUFX4_1210 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_), .Y(adder_bOperand_1_bF_buf0) );
	BUFX4 BUFX4_1211 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .Y(_3675__bF_buf4) );
	BUFX4 BUFX4_1212 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .Y(_3675__bF_buf3) );
	BUFX4 BUFX4_1213 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .Y(_3675__bF_buf2) );
	BUFX4 BUFX4_1214 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .Y(_3675__bF_buf1) );
	BUFX4 BUFX4_1215 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .Y(_3675__bF_buf0) );
	BUFX4 BUFX4_1216 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .Y(_4011__bF_buf3) );
	BUFX4 BUFX4_1217 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .Y(_4011__bF_buf2) );
	BUFX4 BUFX4_1218 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .Y(_4011__bF_buf1) );
	BUFX4 BUFX4_1219 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .Y(_4011__bF_buf0) );
	BUFX4 BUFX4_1220 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_), .Y(divider_divuResult_9_bF_buf5) );
	BUFX4 BUFX4_1221 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_), .Y(divider_divuResult_9_bF_buf4) );
	BUFX4 BUFX4_1222 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_), .Y(divider_divuResult_9_bF_buf3) );
	BUFX4 BUFX4_1223 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_), .Y(divider_divuResult_9_bF_buf2) );
	BUFX4 BUFX4_1224 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_), .Y(divider_divuResult_9_bF_buf1) );
	BUFX4 BUFX4_1225 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_), .Y(divider_divuResult_9_bF_buf0) );
	BUFX4 BUFX4_1226 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .Y(_1517__bF_buf3) );
	BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .Y(_1517__bF_buf2) );
	BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .Y(_1517__bF_buf1) );
	BUFX4 BUFX4_1227 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .Y(_1517__bF_buf0) );
	BUFX4 BUFX4_1228 ( .gnd(gnd), .vdd(vdd), .A(_20629_), .Y(_20629__bF_buf4) );
	BUFX4 BUFX4_1229 ( .gnd(gnd), .vdd(vdd), .A(_20629_), .Y(_20629__bF_buf3) );
	BUFX4 BUFX4_1230 ( .gnd(gnd), .vdd(vdd), .A(_20629_), .Y(_20629__bF_buf2) );
	BUFX4 BUFX4_1231 ( .gnd(gnd), .vdd(vdd), .A(_20629_), .Y(_20629__bF_buf1) );
	BUFX4 BUFX4_1232 ( .gnd(gnd), .vdd(vdd), .A(_20629_), .Y(_20629__bF_buf0) );
	BUFX4 BUFX4_1233 ( .gnd(gnd), .vdd(vdd), .A(_17449_), .Y(_17449__bF_buf4) );
	BUFX4 BUFX4_1234 ( .gnd(gnd), .vdd(vdd), .A(_17449_), .Y(_17449__bF_buf3) );
	BUFX4 BUFX4_1235 ( .gnd(gnd), .vdd(vdd), .A(_17449_), .Y(_17449__bF_buf2) );
	BUFX4 BUFX4_1236 ( .gnd(gnd), .vdd(vdd), .A(_17449_), .Y(_17449__bF_buf1) );
	BUFX4 BUFX4_1237 ( .gnd(gnd), .vdd(vdd), .A(_17449_), .Y(_17449__bF_buf0) );
	BUFX4 BUFX4_1238 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_1746__bF_buf5) );
	BUFX4 BUFX4_1239 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_1746__bF_buf4) );
	BUFX4 BUFX4_1240 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_1746__bF_buf3) );
	BUFX4 BUFX4_1241 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_1746__bF_buf2) );
	BUFX4 BUFX4_1242 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_1746__bF_buf1) );
	BUFX4 BUFX4_1243 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_1746__bF_buf0) );
	BUFX4 BUFX4_1244 ( .gnd(gnd), .vdd(vdd), .A(_17419_), .Y(_17419__bF_buf4) );
	BUFX4 BUFX4_1245 ( .gnd(gnd), .vdd(vdd), .A(_17419_), .Y(_17419__bF_buf3) );
	BUFX4 BUFX4_1246 ( .gnd(gnd), .vdd(vdd), .A(_17419_), .Y(_17419__bF_buf2) );
	BUFX4 BUFX4_1247 ( .gnd(gnd), .vdd(vdd), .A(_17419_), .Y(_17419__bF_buf1) );
	BUFX4 BUFX4_1248 ( .gnd(gnd), .vdd(vdd), .A(_17419_), .Y(_17419__bF_buf0) );
	BUFX4 BUFX4_1249 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_69__bF_buf4) );
	BUFX4 BUFX4_1250 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_69__bF_buf3) );
	BUFX4 BUFX4_1251 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_69__bF_buf2) );
	BUFX4 BUFX4_1252 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_69__bF_buf1) );
	BUFX4 BUFX4_1253 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_69__bF_buf0) );
	BUFX4 BUFX4_1254 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf7) );
	BUFX4 BUFX4_1255 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf6) );
	BUFX4 BUFX4_1256 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf5) );
	BUFX4 BUFX4_1257 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf4) );
	BUFX4 BUFX4_1258 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf3) );
	BUFX4 BUFX4_1259 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf2) );
	BUFX4 BUFX4_1260 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf1) );
	BUFX4 BUFX4_1261 ( .gnd(gnd), .vdd(vdd), .A(_20557_), .Y(_20557__bF_buf0) );
	BUFX4 BUFX4_1262 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf6) );
	BUFX4 BUFX4_1263 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf5) );
	BUFX4 BUFX4_1264 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf4) );
	BUFX4 BUFX4_1265 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf3) );
	BUFX4 BUFX4_1266 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf2) );
	BUFX4 BUFX4_1267 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf1) );
	BUFX4 BUFX4_1268 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_), .Y(divider_divuResult_4_bF_buf0) );
	BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_), .Y(aOperand_frameOut_25_bF_buf3) );
	BUFX4 BUFX4_1269 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_), .Y(aOperand_frameOut_25_bF_buf2) );
	BUFX4 BUFX4_1270 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_), .Y(aOperand_frameOut_25_bF_buf1) );
	BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_), .Y(aOperand_frameOut_25_bF_buf0) );
	BUFX4 BUFX4_1271 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf7) );
	BUFX4 BUFX4_1272 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf6) );
	BUFX4 BUFX4_1273 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf5) );
	BUFX4 BUFX4_1274 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf4) );
	BUFX4 BUFX4_1275 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf3) );
	BUFX4 BUFX4_1276 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf2) );
	BUFX4 BUFX4_1277 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf1) );
	BUFX4 BUFX4_1278 ( .gnd(gnd), .vdd(vdd), .A(_20425_), .Y(_20425__bF_buf0) );
	BUFX4 BUFX4_1279 ( .gnd(gnd), .vdd(vdd), .A(_20624_), .Y(_20624__bF_buf4) );
	BUFX4 BUFX4_1280 ( .gnd(gnd), .vdd(vdd), .A(_20624_), .Y(_20624__bF_buf3) );
	BUFX4 BUFX4_1281 ( .gnd(gnd), .vdd(vdd), .A(_20624_), .Y(_20624__bF_buf2) );
	BUFX4 BUFX4_1282 ( .gnd(gnd), .vdd(vdd), .A(_20624_), .Y(_20624__bF_buf1) );
	BUFX4 BUFX4_1283 ( .gnd(gnd), .vdd(vdd), .A(_20624_), .Y(_20624__bF_buf0) );
	BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_), .Y(aOperand_frameOut_20_bF_buf4) );
	BUFX4 BUFX4_1284 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_), .Y(aOperand_frameOut_20_bF_buf3) );
	BUFX4 BUFX4_1285 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_), .Y(aOperand_frameOut_20_bF_buf2) );
	BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_), .Y(aOperand_frameOut_20_bF_buf1) );
	BUFX4 BUFX4_1286 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_), .Y(aOperand_frameOut_20_bF_buf0) );
	BUFX4 BUFX4_1287 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .Y(_4937__bF_buf5) );
	BUFX4 BUFX4_1288 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .Y(_4937__bF_buf4) );
	BUFX4 BUFX4_1289 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .Y(_4937__bF_buf3) );
	BUFX4 BUFX4_1290 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .Y(_4937__bF_buf2) );
	BUFX4 BUFX4_1291 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .Y(_4937__bF_buf1) );
	BUFX4 BUFX4_1292 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .Y(_4937__bF_buf0) );
	BUFX4 BUFX4_1293 ( .gnd(gnd), .vdd(vdd), .A(_4504_), .Y(_4504__bF_buf4) );
	BUFX4 BUFX4_1294 ( .gnd(gnd), .vdd(vdd), .A(_4504_), .Y(_4504__bF_buf3) );
	BUFX4 BUFX4_1295 ( .gnd(gnd), .vdd(vdd), .A(_4504_), .Y(_4504__bF_buf2) );
	BUFX4 BUFX4_1296 ( .gnd(gnd), .vdd(vdd), .A(_4504_), .Y(_4504__bF_buf1) );
	BUFX4 BUFX4_1297 ( .gnd(gnd), .vdd(vdd), .A(_4504_), .Y(_4504__bF_buf0) );
	BUFX4 BUFX4_1298 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf7) );
	BUFX4 BUFX4_1299 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf6) );
	BUFX4 BUFX4_1300 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf5) );
	BUFX4 BUFX4_1301 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf4) );
	BUFX4 BUFX4_1302 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf3) );
	BUFX4 BUFX4_1303 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf2) );
	BUFX4 BUFX4_1304 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf1) );
	BUFX4 BUFX4_1305 ( .gnd(gnd), .vdd(vdd), .A(_19769_), .Y(_19769__bF_buf0) );
	BUFX4 BUFX4_1306 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf7) );
	BUFX4 BUFX4_1307 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf6) );
	BUFX4 BUFX4_1308 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf5) );
	BUFX4 BUFX4_1309 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf4) );
	BUFX4 BUFX4_1310 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf3) );
	BUFX4 BUFX4_1311 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf2) );
	BUFX4 BUFX4_1312 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf1) );
	BUFX4 BUFX4_1313 ( .gnd(gnd), .vdd(vdd), .A(_19396_), .Y(_19396__bF_buf0) );
	BUFX4 BUFX4_1314 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf7) );
	BUFX4 BUFX4_1315 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf6) );
	BUFX4 BUFX4_1316 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf5) );
	BUFX4 BUFX4_1317 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf4) );
	BUFX4 BUFX4_1318 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf3) );
	BUFX4 BUFX4_1319 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf2) );
	BUFX4 BUFX4_1320 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf1) );
	BUFX4 BUFX4_1321 ( .gnd(gnd), .vdd(vdd), .A(_19968_), .Y(_19968__bF_buf0) );
	BUFX4 BUFX4_1322 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_), .Y(aOperand_frameOut_18_bF_buf4) );
	BUFX4 BUFX4_1323 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_), .Y(aOperand_frameOut_18_bF_buf3) );
	BUFX4 BUFX4_1324 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_), .Y(aOperand_frameOut_18_bF_buf2) );
	BUFX4 BUFX4_1325 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_), .Y(aOperand_frameOut_18_bF_buf1) );
	BUFX4 BUFX4_1326 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_), .Y(aOperand_frameOut_18_bF_buf0) );
	BUFX4 BUFX4_1327 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .Y(_1505__bF_buf4) );
	BUFX4 BUFX4_1328 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .Y(_1505__bF_buf3) );
	BUFX4 BUFX4_1329 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .Y(_1505__bF_buf2) );
	BUFX4 BUFX4_1330 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .Y(_1505__bF_buf1) );
	BUFX4 BUFX4_1331 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .Y(_1505__bF_buf0) );
	BUFX4 BUFX4_1332 ( .gnd(gnd), .vdd(vdd), .A(_20617_), .Y(_20617__bF_buf4) );
	BUFX4 BUFX4_1333 ( .gnd(gnd), .vdd(vdd), .A(_20617_), .Y(_20617__bF_buf3) );
	BUFX4 BUFX4_1334 ( .gnd(gnd), .vdd(vdd), .A(_20617_), .Y(_20617__bF_buf2) );
	BUFX4 BUFX4_1335 ( .gnd(gnd), .vdd(vdd), .A(_20617_), .Y(_20617__bF_buf1) );
	BUFX4 BUFX4_1336 ( .gnd(gnd), .vdd(vdd), .A(_20617_), .Y(_20617__bF_buf0) );
	BUFX4 BUFX4_1337 ( .gnd(gnd), .vdd(vdd), .A(_17467_), .Y(_17467__bF_buf4) );
	BUFX4 BUFX4_1338 ( .gnd(gnd), .vdd(vdd), .A(_17467_), .Y(_17467__bF_buf3) );
	BUFX4 BUFX4_1339 ( .gnd(gnd), .vdd(vdd), .A(_17467_), .Y(_17467__bF_buf2) );
	BUFX4 BUFX4_1340 ( .gnd(gnd), .vdd(vdd), .A(_17467_), .Y(_17467__bF_buf1) );
	BUFX4 BUFX4_1341 ( .gnd(gnd), .vdd(vdd), .A(_17467_), .Y(_17467__bF_buf0) );
	BUFX4 BUFX4_1342 ( .gnd(gnd), .vdd(vdd), .A(_17407_), .Y(_17407__bF_buf4) );
	BUFX4 BUFX4_1343 ( .gnd(gnd), .vdd(vdd), .A(_17407_), .Y(_17407__bF_buf3) );
	BUFX4 BUFX4_1344 ( .gnd(gnd), .vdd(vdd), .A(_17407_), .Y(_17407__bF_buf2) );
	BUFX4 BUFX4_1345 ( .gnd(gnd), .vdd(vdd), .A(_17407_), .Y(_17407__bF_buf1) );
	BUFX4 BUFX4_1346 ( .gnd(gnd), .vdd(vdd), .A(_17407_), .Y(_17407__bF_buf0) );
	BUFX4 BUFX4_1347 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf3) );
	BUFX4 BUFX4_1348 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf2) );
	BUFX4 BUFX4_1349 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf1) );
	BUFX4 BUFX4_1350 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf0) );
	BUFX4 BUFX4_1351 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_), .Y(divider_absoluteValue_B_flipSign_result_23_bF_buf3) );
	BUFX4 BUFX4_1352 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_), .Y(divider_absoluteValue_B_flipSign_result_23_bF_buf2) );
	BUFX4 BUFX4_1353 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_), .Y(divider_absoluteValue_B_flipSign_result_23_bF_buf1) );
	BUFX4 BUFX4_1354 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_), .Y(divider_absoluteValue_B_flipSign_result_23_bF_buf0) );
	BUFX4 BUFX4_1355 ( .gnd(gnd), .vdd(vdd), .A(_20575_), .Y(_20575__bF_buf4) );
	BUFX4 BUFX4_1356 ( .gnd(gnd), .vdd(vdd), .A(_20575_), .Y(_20575__bF_buf3) );
	BUFX4 BUFX4_1357 ( .gnd(gnd), .vdd(vdd), .A(_20575_), .Y(_20575__bF_buf2) );
	BUFX4 BUFX4_1358 ( .gnd(gnd), .vdd(vdd), .A(_20575_), .Y(_20575__bF_buf1) );
	BUFX4 BUFX4_1359 ( .gnd(gnd), .vdd(vdd), .A(_20575_), .Y(_20575__bF_buf0) );
	BUFX4 BUFX4_1360 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf7) );
	BUFX4 BUFX4_1361 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf6) );
	BUFX4 BUFX4_1362 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf5) );
	BUFX4 BUFX4_1363 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf4) );
	BUFX4 BUFX4_1364 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf3) );
	BUFX4 BUFX4_1365 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf2) );
	BUFX4 BUFX4_1366 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf1) );
	BUFX4 BUFX4_1367 ( .gnd(gnd), .vdd(vdd), .A(_19602_), .Y(_19602__bF_buf0) );
	BUFX4 BUFX4_1368 ( .gnd(gnd), .vdd(vdd), .A(_11712_), .Y(_11712__bF_buf4) );
	BUFX4 BUFX4_1369 ( .gnd(gnd), .vdd(vdd), .A(_11712_), .Y(_11712__bF_buf3) );
	BUFX4 BUFX4_1370 ( .gnd(gnd), .vdd(vdd), .A(_11712_), .Y(_11712__bF_buf2) );
	BUFX4 BUFX4_1371 ( .gnd(gnd), .vdd(vdd), .A(_11712_), .Y(_11712__bF_buf1) );
	BUFX4 BUFX4_1372 ( .gnd(gnd), .vdd(vdd), .A(_11712_), .Y(_11712__bF_buf0) );
	BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_), .Y(adder_bOperand_21_bF_buf3) );
	BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_), .Y(adder_bOperand_21_bF_buf2) );
	BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_), .Y(adder_bOperand_21_bF_buf1) );
	BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_), .Y(adder_bOperand_21_bF_buf0) );
	BUFX4 BUFX4_1373 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_), .Y(aOperand_frameOut_13_bF_buf4) );
	BUFX4 BUFX4_1374 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_), .Y(aOperand_frameOut_13_bF_buf3) );
	BUFX4 BUFX4_1375 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_), .Y(aOperand_frameOut_13_bF_buf2) );
	BUFX4 BUFX4_1376 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_), .Y(aOperand_frameOut_13_bF_buf1) );
	BUFX4 BUFX4_1377 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_), .Y(aOperand_frameOut_13_bF_buf0) );
	BUFX4 BUFX4_1378 ( .gnd(gnd), .vdd(vdd), .A(_11971_), .Y(_11971__bF_buf3) );
	BUFX4 BUFX4_1379 ( .gnd(gnd), .vdd(vdd), .A(_11971_), .Y(_11971__bF_buf2) );
	BUFX4 BUFX4_1380 ( .gnd(gnd), .vdd(vdd), .A(_11971_), .Y(_11971__bF_buf1) );
	BUFX4 BUFX4_1381 ( .gnd(gnd), .vdd(vdd), .A(_11971_), .Y(_11971__bF_buf0) );
	BUFX4 BUFX4_1382 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_), .Y(aOperand_frameOut_8_bF_buf4) );
	BUFX4 BUFX4_1383 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_), .Y(aOperand_frameOut_8_bF_buf3) );
	BUFX4 BUFX4_1384 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_), .Y(aOperand_frameOut_8_bF_buf2) );
	BUFX4 BUFX4_1385 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_), .Y(aOperand_frameOut_8_bF_buf1) );
	BUFX4 BUFX4_1386 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_), .Y(aOperand_frameOut_8_bF_buf0) );
	BUFX4 BUFX4_1387 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .Y(_1560__bF_buf3) );
	BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .Y(_1560__bF_buf2) );
	BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .Y(_1560__bF_buf1) );
	BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .Y(_1560__bF_buf0) );
	BUFX4 BUFX4_1388 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_), .Y(reg_dataIn_26_bF_buf4) );
	BUFX4 BUFX4_1389 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_), .Y(reg_dataIn_26_bF_buf3) );
	BUFX4 BUFX4_1390 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_), .Y(reg_dataIn_26_bF_buf2) );
	BUFX4 BUFX4_1391 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_), .Y(reg_dataIn_26_bF_buf1) );
	BUFX4 BUFX4_1392 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_), .Y(reg_dataIn_26_bF_buf0) );
	BUFX4 BUFX4_1393 ( .gnd(gnd), .vdd(vdd), .A(_17462_), .Y(_17462__bF_buf4) );
	BUFX4 BUFX4_1394 ( .gnd(gnd), .vdd(vdd), .A(_17462_), .Y(_17462__bF_buf3) );
	BUFX4 BUFX4_1395 ( .gnd(gnd), .vdd(vdd), .A(_17462_), .Y(_17462__bF_buf2) );
	BUFX4 BUFX4_1396 ( .gnd(gnd), .vdd(vdd), .A(_17462_), .Y(_17462__bF_buf1) );
	BUFX4 BUFX4_1397 ( .gnd(gnd), .vdd(vdd), .A(_17462_), .Y(_17462__bF_buf0) );
	BUFX4 BUFX4_1398 ( .gnd(gnd), .vdd(vdd), .A(_17432_), .Y(_17432__bF_buf4) );
	BUFX4 BUFX4_1399 ( .gnd(gnd), .vdd(vdd), .A(_17432_), .Y(_17432__bF_buf3) );
	BUFX4 BUFX4_1400 ( .gnd(gnd), .vdd(vdd), .A(_17432_), .Y(_17432__bF_buf2) );
	BUFX4 BUFX4_1401 ( .gnd(gnd), .vdd(vdd), .A(_17432_), .Y(_17432__bF_buf1) );
	BUFX4 BUFX4_1402 ( .gnd(gnd), .vdd(vdd), .A(_17432_), .Y(_17432__bF_buf0) );
	BUFX4 BUFX4_1403 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_82__bF_buf4) );
	BUFX4 BUFX4_1404 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_82__bF_buf3) );
	BUFX4 BUFX4_1405 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_82__bF_buf2) );
	BUFX4 BUFX4_1406 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_82__bF_buf1) );
	BUFX4 BUFX4_1407 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_82__bF_buf0) );
	BUFX4 BUFX4_1408 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .Y(_5886__bF_buf3) );
	BUFX4 BUFX4_1409 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .Y(_5886__bF_buf2) );
	BUFX4 BUFX4_1410 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .Y(_5886__bF_buf1) );
	BUFX4 BUFX4_1411 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .Y(_5886__bF_buf0) );
	BUFX4 BUFX4_1412 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_), .Y(aOperand_frameOut_3_bF_buf4) );
	BUFX4 BUFX4_1413 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_), .Y(aOperand_frameOut_3_bF_buf3) );
	BUFX4 BUFX4_1414 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_), .Y(aOperand_frameOut_3_bF_buf2) );
	BUFX4 BUFX4_1415 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_), .Y(aOperand_frameOut_3_bF_buf1) );
	BUFX4 BUFX4_1416 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_), .Y(aOperand_frameOut_3_bF_buf0) );
	BUFX4 BUFX4_1417 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_), .Y(reg_dataIn_21_bF_buf4) );
	BUFX4 BUFX4_1418 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_), .Y(reg_dataIn_21_bF_buf3) );
	BUFX4 BUFX4_1419 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_), .Y(reg_dataIn_21_bF_buf2) );
	BUFX4 BUFX4_1420 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_), .Y(reg_dataIn_21_bF_buf1) );
	BUFX4 BUFX4_1421 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_), .Y(reg_dataIn_21_bF_buf0) );
	BUFX4 BUFX4_1422 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_), .Y(divider_divuResult_24_bF_buf3) );
	BUFX4 BUFX4_1423 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_), .Y(divider_divuResult_24_bF_buf2) );
	BUFX4 BUFX4_1424 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_), .Y(divider_divuResult_24_bF_buf1) );
	BUFX4 BUFX4_1425 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_), .Y(divider_divuResult_24_bF_buf0) );
	BUFX4 BUFX4_1426 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_), .Y(adder_bOperand_19_bF_buf3) );
	BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_), .Y(adder_bOperand_19_bF_buf2) );
	BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_), .Y(adder_bOperand_19_bF_buf1) );
	BUFX4 BUFX4_1427 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_), .Y(adder_bOperand_19_bF_buf0) );
	BUFX4 BUFX4_1428 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .Y(_2887__bF_buf4) );
	BUFX4 BUFX4_1429 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .Y(_2887__bF_buf3) );
	BUFX4 BUFX4_1430 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .Y(_2887__bF_buf2) );
	BUFX4 BUFX4_1431 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .Y(_2887__bF_buf1) );
	BUFX4 BUFX4_1432 ( .gnd(gnd), .vdd(vdd), .A(_2887_), .Y(_2887__bF_buf0) );
	BUFX4 BUFX4_1433 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .Y(_2255__bF_buf4) );
	BUFX4 BUFX4_1434 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .Y(_2255__bF_buf3) );
	BUFX4 BUFX4_1435 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .Y(_2255__bF_buf2) );
	BUFX4 BUFX4_1436 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .Y(_2255__bF_buf1) );
	BUFX4 BUFX4_1437 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .Y(_2255__bF_buf0) );
	BUFX4 BUFX4_1438 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_), .Y(reg_dataIn_9_bF_buf4) );
	BUFX4 BUFX4_1439 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_), .Y(reg_dataIn_9_bF_buf3) );
	BUFX4 BUFX4_1440 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_), .Y(reg_dataIn_9_bF_buf2) );
	BUFX4 BUFX4_1441 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_), .Y(reg_dataIn_9_bF_buf1) );
	BUFX4 BUFX4_1442 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_), .Y(reg_dataIn_9_bF_buf0) );
	BUFX4 BUFX4_1443 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .Y(_1757__bF_buf3) );
	BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .Y(_1757__bF_buf2) );
	BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .Y(_1757__bF_buf1) );
	BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .Y(_1757__bF_buf0) );
	BUFX4 BUFX4_1444 ( .gnd(gnd), .vdd(vdd), .A(_20598_), .Y(_20598__bF_buf4) );
	BUFX4 BUFX4_1445 ( .gnd(gnd), .vdd(vdd), .A(_20598_), .Y(_20598__bF_buf3) );
	BUFX4 BUFX4_1446 ( .gnd(gnd), .vdd(vdd), .A(_20598_), .Y(_20598__bF_buf2) );
	BUFX4 BUFX4_1447 ( .gnd(gnd), .vdd(vdd), .A(_20598_), .Y(_20598__bF_buf1) );
	BUFX4 BUFX4_1448 ( .gnd(gnd), .vdd(vdd), .A(_20598_), .Y(_20598__bF_buf0) );
	BUFX4 BUFX4_1449 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_), .Y(divider_absoluteValue_B_flipSign_result_16_bF_buf5) );
	BUFX4 BUFX4_1450 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_), .Y(divider_absoluteValue_B_flipSign_result_16_bF_buf4) );
	BUFX4 BUFX4_1451 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_), .Y(divider_absoluteValue_B_flipSign_result_16_bF_buf3) );
	BUFX4 BUFX4_1452 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_), .Y(divider_absoluteValue_B_flipSign_result_16_bF_buf2) );
	BUFX4 BUFX4_1453 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_), .Y(divider_absoluteValue_B_flipSign_result_16_bF_buf1) );
	BUFX4 BUFX4_1454 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_), .Y(divider_absoluteValue_B_flipSign_result_16_bF_buf0) );
	BUFX4 BUFX4_1455 ( .gnd(gnd), .vdd(vdd), .A(_20568_), .Y(_20568__bF_buf4) );
	BUFX4 BUFX4_1456 ( .gnd(gnd), .vdd(vdd), .A(_20568_), .Y(_20568__bF_buf3) );
	BUFX4 BUFX4_1457 ( .gnd(gnd), .vdd(vdd), .A(_20568_), .Y(_20568__bF_buf2) );
	BUFX4 BUFX4_1458 ( .gnd(gnd), .vdd(vdd), .A(_20568_), .Y(_20568__bF_buf1) );
	BUFX4 BUFX4_1459 ( .gnd(gnd), .vdd(vdd), .A(_20568_), .Y(_20568__bF_buf0) );
	BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_), .Y(adder_bOperand_14_bF_buf3) );
	BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_), .Y(adder_bOperand_14_bF_buf2) );
	BUFX4 BUFX4_1460 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_), .Y(adder_bOperand_14_bF_buf1) );
	BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_), .Y(adder_bOperand_14_bF_buf0) );
	BUFX4 BUFX4_1461 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_), .Y(reg_dataIn_4_bF_buf4) );
	BUFX4 BUFX4_1462 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_), .Y(reg_dataIn_4_bF_buf3) );
	BUFX4 BUFX4_1463 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_), .Y(reg_dataIn_4_bF_buf2) );
	BUFX4 BUFX4_1464 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_), .Y(reg_dataIn_4_bF_buf1) );
	BUFX4 BUFX4_1465 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_), .Y(reg_dataIn_4_bF_buf0) );
	BUFX4 BUFX4_1466 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_), .Y(reg_dataIn_19_bF_buf4) );
	BUFX4 BUFX4_1467 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_), .Y(reg_dataIn_19_bF_buf3) );
	BUFX4 BUFX4_1468 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_), .Y(reg_dataIn_19_bF_buf2) );
	BUFX4 BUFX4_1469 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_), .Y(reg_dataIn_19_bF_buf1) );
	BUFX4 BUFX4_1470 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_), .Y(reg_dataIn_19_bF_buf0) );
	BUFX4 BUFX4_1471 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf6) );
	BUFX4 BUFX4_1472 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf5) );
	BUFX4 BUFX4_1473 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf4) );
	BUFX4 BUFX4_1474 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf3) );
	BUFX4 BUFX4_1475 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf2) );
	BUFX4 BUFX4_1476 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf1) );
	BUFX4 BUFX4_1477 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_), .Y(divider_absoluteValue_B_flipSign_result_9_bF_buf0) );
	BUFX4 BUFX4_1478 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9913__bF_buf5) );
	BUFX4 BUFX4_1479 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9913__bF_buf4) );
	BUFX4 BUFX4_1480 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9913__bF_buf3) );
	BUFX4 BUFX4_1481 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9913__bF_buf2) );
	BUFX4 BUFX4_1482 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9913__bF_buf1) );
	BUFX4 BUFX4_1483 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .Y(_9913__bF_buf0) );
	BUFX4 BUFX4_1484 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_), .Y(divider_absoluteValue_B_flipSign_result_11_bF_buf5) );
	BUFX4 BUFX4_1485 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_), .Y(divider_absoluteValue_B_flipSign_result_11_bF_buf4) );
	BUFX4 BUFX4_1486 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_), .Y(divider_absoluteValue_B_flipSign_result_11_bF_buf3) );
	BUFX4 BUFX4_1487 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_), .Y(divider_absoluteValue_B_flipSign_result_11_bF_buf2) );
	BUFX4 BUFX4_1488 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_), .Y(divider_absoluteValue_B_flipSign_result_11_bF_buf1) );
	BUFX4 BUFX4_1489 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_), .Y(divider_absoluteValue_B_flipSign_result_11_bF_buf0) );
	BUFX4 BUFX4_1490 ( .gnd(gnd), .vdd(vdd), .A(_17383_), .Y(_17383__bF_buf4) );
	BUFX4 BUFX4_1491 ( .gnd(gnd), .vdd(vdd), .A(_17383_), .Y(_17383__bF_buf3) );
	BUFX4 BUFX4_1492 ( .gnd(gnd), .vdd(vdd), .A(_17383_), .Y(_17383__bF_buf2) );
	BUFX4 BUFX4_1493 ( .gnd(gnd), .vdd(vdd), .A(_17383_), .Y(_17383__bF_buf1) );
	BUFX4 BUFX4_1494 ( .gnd(gnd), .vdd(vdd), .A(_17383_), .Y(_17383__bF_buf0) );
	BUFX4 BUFX4_1495 ( .gnd(gnd), .vdd(vdd), .A(_17022_), .Y(_17022__bF_buf3) );
	BUFX4 BUFX4_1496 ( .gnd(gnd), .vdd(vdd), .A(_17022_), .Y(_17022__bF_buf2) );
	BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_17022_), .Y(_17022__bF_buf1) );
	BUFX4 BUFX4_1497 ( .gnd(gnd), .vdd(vdd), .A(_17022_), .Y(_17022__bF_buf0) );
	BUFX4 BUFX4_1498 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_), .Y(reg_dataIn_14_bF_buf4) );
	BUFX4 BUFX4_1499 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_), .Y(reg_dataIn_14_bF_buf3) );
	BUFX4 BUFX4_1500 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_), .Y(reg_dataIn_14_bF_buf2) );
	BUFX4 BUFX4_1501 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_), .Y(reg_dataIn_14_bF_buf1) );
	BUFX4 BUFX4_1502 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_), .Y(reg_dataIn_14_bF_buf0) );
	BUFX4 BUFX4_1503 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_17_), .Y(divider_divuResult_17_bF_buf3) );
	BUFX4 BUFX4_1504 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_17_), .Y(divider_divuResult_17_bF_buf2) );
	BUFX4 BUFX4_1505 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_17_), .Y(divider_divuResult_17_bF_buf1) );
	BUFX4 BUFX4_1506 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_17_), .Y(divider_divuResult_17_bF_buf0) );
	BUFX4 BUFX4_1507 ( .gnd(gnd), .vdd(vdd), .A(_20630_), .Y(_20630__bF_buf4) );
	BUFX4 BUFX4_1508 ( .gnd(gnd), .vdd(vdd), .A(_20630_), .Y(_20630__bF_buf3) );
	BUFX4 BUFX4_1509 ( .gnd(gnd), .vdd(vdd), .A(_20630_), .Y(_20630__bF_buf2) );
	BUFX4 BUFX4_1510 ( .gnd(gnd), .vdd(vdd), .A(_20630_), .Y(_20630__bF_buf1) );
	BUFX4 BUFX4_1511 ( .gnd(gnd), .vdd(vdd), .A(_20630_), .Y(_20630__bF_buf0) );
	BUFX4 BUFX4_1512 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf6) );
	BUFX4 BUFX4_1513 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf5) );
	BUFX4 BUFX4_1514 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf4) );
	BUFX4 BUFX4_1515 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf3) );
	BUFX4 BUFX4_1516 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf2) );
	BUFX4 BUFX4_1517 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf1) );
	BUFX4 BUFX4_1518 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_), .Y(divider_absoluteValue_B_flipSign_result_4_bF_buf0) );
	BUFX4 BUFX4_1519 ( .gnd(gnd), .vdd(vdd), .A(_17450_), .Y(_17450__bF_buf4) );
	BUFX4 BUFX4_1520 ( .gnd(gnd), .vdd(vdd), .A(_17450_), .Y(_17450__bF_buf3) );
	BUFX4 BUFX4_1521 ( .gnd(gnd), .vdd(vdd), .A(_17450_), .Y(_17450__bF_buf2) );
	BUFX4 BUFX4_1522 ( .gnd(gnd), .vdd(vdd), .A(_17450_), .Y(_17450__bF_buf1) );
	BUFX4 BUFX4_1523 ( .gnd(gnd), .vdd(vdd), .A(_17450_), .Y(_17450__bF_buf0) );
	BUFX4 BUFX4_1524 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .Y(_6342__bF_buf4) );
	BUFX4 BUFX4_1525 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .Y(_6342__bF_buf3) );
	BUFX4 BUFX4_1526 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .Y(_6342__bF_buf2) );
	BUFX4 BUFX4_1527 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .Y(_6342__bF_buf1) );
	BUFX4 BUFX4_1528 ( .gnd(gnd), .vdd(vdd), .A(_6342_), .Y(_6342__bF_buf0) );
	BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_), .Y(adder_bOperand_5_bF_buf4) );
	BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_), .Y(adder_bOperand_5_bF_buf3) );
	BUFX4 BUFX4_1529 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_), .Y(adder_bOperand_5_bF_buf2) );
	BUFX4 BUFX4_1530 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_), .Y(adder_bOperand_5_bF_buf1) );
	BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_), .Y(adder_bOperand_5_bF_buf0) );
	BUFX4 BUFX4_1531 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf6) );
	BUFX4 BUFX4_1532 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf5) );
	BUFX4 BUFX4_1533 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf4) );
	BUFX4 BUFX4_1534 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf3) );
	BUFX4 BUFX4_1535 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf2) );
	BUFX4 BUFX4_1536 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf1) );
	BUFX4 BUFX4_1537 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_), .Y(divider_divuResult_12_bF_buf0) );
	BUFX4 BUFX4_1538 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf6) );
	BUFX4 BUFX4_1539 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf5) );
	BUFX4 BUFX4_1540 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf4) );
	BUFX4 BUFX4_1541 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf3) );
	BUFX4 BUFX4_1542 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf2) );
	BUFX4 BUFX4_1543 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf1) );
	BUFX4 BUFX4_1544 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .Y(_4714__bF_buf0) );
	BUFX4 BUFX4_1545 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf6) );
	BUFX4 BUFX4_1546 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf5) );
	BUFX4 BUFX4_1547 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf4) );
	BUFX4 BUFX4_1548 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf3) );
	BUFX4 BUFX4_1549 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf2) );
	BUFX4 BUFX4_1550 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf1) );
	BUFX4 BUFX4_1551 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_), .Y(adder_bOperand_0_bF_buf0) );
	BUFX4 BUFX4_1552 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .Y(_4010__bF_buf4) );
	BUFX4 BUFX4_1553 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .Y(_4010__bF_buf3) );
	BUFX4 BUFX4_1554 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .Y(_4010__bF_buf2) );
	BUFX4 BUFX4_1555 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .Y(_4010__bF_buf1) );
	BUFX4 BUFX4_1556 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .Y(_4010__bF_buf0) );
	BUFX4 BUFX4_1557 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf6) );
	BUFX4 BUFX4_1558 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf5) );
	BUFX4 BUFX4_1559 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf4) );
	BUFX4 BUFX4_1560 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf3) );
	BUFX4 BUFX4_1561 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf2) );
	BUFX4 BUFX4_1562 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf1) );
	BUFX4 BUFX4_1563 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_), .Y(divider_divuResult_8_bF_buf0) );
	BUFX4 BUFX4_1564 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .Y(_2917__bF_buf4) );
	BUFX4 BUFX4_1565 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .Y(_2917__bF_buf3) );
	BUFX4 BUFX4_1566 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .Y(_2917__bF_buf2) );
	BUFX4 BUFX4_1567 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .Y(_2917__bF_buf1) );
	BUFX4 BUFX4_1568 ( .gnd(gnd), .vdd(vdd), .A(_2917_), .Y(_2917__bF_buf0) );
	BUFX4 BUFX4_1569 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .Y(_12353__bF_buf3) );
	BUFX4 BUFX4_1570 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .Y(_12353__bF_buf2) );
	BUFX4 BUFX4_1571 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .Y(_12353__bF_buf1) );
	BUFX4 BUFX4_1572 ( .gnd(gnd), .vdd(vdd), .A(_12353_), .Y(_12353__bF_buf0) );
	BUFX4 BUFX4_1573 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .Y(_11054__bF_buf4) );
	BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .Y(_11054__bF_buf3) );
	BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .Y(_11054__bF_buf2) );
	BUFX4 BUFX4_1574 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .Y(_11054__bF_buf1) );
	BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .Y(_11054__bF_buf0) );
	BUFX4 BUFX4_1575 ( .gnd(gnd), .vdd(vdd), .A(_8697_), .Y(_8697__bF_buf3) );
	BUFX4 BUFX4_1576 ( .gnd(gnd), .vdd(vdd), .A(_8697_), .Y(_8697__bF_buf2) );
	BUFX4 BUFX4_1577 ( .gnd(gnd), .vdd(vdd), .A(_8697_), .Y(_8697__bF_buf1) );
	BUFX4 BUFX4_1578 ( .gnd(gnd), .vdd(vdd), .A(_8697_), .Y(_8697__bF_buf0) );
	BUFX4 BUFX4_1579 ( .gnd(gnd), .vdd(vdd), .A(_17418_), .Y(_17418__bF_buf4) );
	BUFX4 BUFX4_1580 ( .gnd(gnd), .vdd(vdd), .A(_17418_), .Y(_17418__bF_buf3) );
	BUFX4 BUFX4_1581 ( .gnd(gnd), .vdd(vdd), .A(_17418_), .Y(_17418__bF_buf2) );
	BUFX4 BUFX4_1582 ( .gnd(gnd), .vdd(vdd), .A(_17418_), .Y(_17418__bF_buf1) );
	BUFX4 BUFX4_1583 ( .gnd(gnd), .vdd(vdd), .A(_17418_), .Y(_17418__bF_buf0) );
	BUFX4 BUFX4_1584 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf4) );
	BUFX4 BUFX4_1585 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf3) );
	BUFX4 BUFX4_1586 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf2) );
	BUFX4 BUFX4_1587 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf1) );
	BUFX4 BUFX4_1588 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf0) );
	BUFX4 BUFX4_1589 ( .gnd(gnd), .vdd(vdd), .A(_20586_), .Y(_20586__bF_buf4) );
	BUFX4 BUFX4_1590 ( .gnd(gnd), .vdd(vdd), .A(_20586_), .Y(_20586__bF_buf3) );
	BUFX4 BUFX4_1591 ( .gnd(gnd), .vdd(vdd), .A(_20586_), .Y(_20586__bF_buf2) );
	BUFX4 BUFX4_1592 ( .gnd(gnd), .vdd(vdd), .A(_20586_), .Y(_20586__bF_buf1) );
	BUFX4 BUFX4_1593 ( .gnd(gnd), .vdd(vdd), .A(_20586_), .Y(_20586__bF_buf0) );
	BUFX4 BUFX4_1594 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .Y(_17376__bF_buf5) );
	BUFX4 BUFX4_1595 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .Y(_17376__bF_buf4) );
	BUFX4 BUFX4_1596 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .Y(_17376__bF_buf3) );
	BUFX4 BUFX4_1597 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .Y(_17376__bF_buf2) );
	BUFX4 BUFX4_1598 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .Y(_17376__bF_buf1) );
	BUFX4 BUFX4_1599 ( .gnd(gnd), .vdd(vdd), .A(_17376_), .Y(_17376__bF_buf0) );
	BUFX4 BUFX4_1600 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf7) );
	BUFX4 BUFX4_1601 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf6) );
	BUFX4 BUFX4_1602 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf5) );
	BUFX4 BUFX4_1603 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf4) );
	BUFX4 BUFX4_1604 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf3) );
	BUFX4 BUFX4_1605 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf2) );
	BUFX4 BUFX4_1606 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf1) );
	BUFX4 BUFX4_1607 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_), .Y(divider_divuResult_3_bF_buf0) );
	BUFX4 BUFX4_1608 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .Y(_1944__bF_buf4) );
	BUFX4 BUFX4_1609 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .Y(_1944__bF_buf3) );
	BUFX4 BUFX4_1610 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .Y(_1944__bF_buf2) );
	BUFX4 BUFX4_1611 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .Y(_1944__bF_buf1) );
	BUFX4 BUFX4_1612 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .Y(_1944__bF_buf0) );
	BUFX4 BUFX4_1613 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_), .Y(aOperand_frameOut_24_bF_buf3) );
	BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_), .Y(aOperand_frameOut_24_bF_buf2) );
	BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_), .Y(aOperand_frameOut_24_bF_buf1) );
	BUFX4 BUFX4_1614 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_), .Y(aOperand_frameOut_24_bF_buf0) );
	BUFX4 BUFX4_1615 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .Y(_5499__bF_buf3) );
	BUFX4 BUFX4_1616 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .Y(_5499__bF_buf2) );
	BUFX4 BUFX4_1617 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .Y(_5499__bF_buf1) );
	BUFX4 BUFX4_1618 ( .gnd(gnd), .vdd(vdd), .A(_5499_), .Y(_5499__bF_buf0) );
	BUFX4 BUFX4_1619 ( .gnd(gnd), .vdd(vdd), .A(_17443_), .Y(_17443__bF_buf4) );
	BUFX4 BUFX4_1620 ( .gnd(gnd), .vdd(vdd), .A(_17443_), .Y(_17443__bF_buf3) );
	BUFX4 BUFX4_1621 ( .gnd(gnd), .vdd(vdd), .A(_17443_), .Y(_17443__bF_buf2) );
	BUFX4 BUFX4_1622 ( .gnd(gnd), .vdd(vdd), .A(_17443_), .Y(_17443__bF_buf1) );
	BUFX4 BUFX4_1623 ( .gnd(gnd), .vdd(vdd), .A(_17443_), .Y(_17443__bF_buf0) );
	BUFX4 BUFX4_1624 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf7) );
	BUFX4 BUFX4_1625 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf6) );
	BUFX4 BUFX4_1626 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf5) );
	BUFX4 BUFX4_1627 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf4) );
	BUFX4 BUFX4_1628 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf3) );
	BUFX4 BUFX4_1629 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf2) );
	BUFX4 BUFX4_1630 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf1) );
	BUFX4 BUFX4_1631 ( .gnd(gnd), .vdd(vdd), .A(_17413_), .Y(_17413__bF_buf0) );
	BUFX4 BUFX4_1632 ( .gnd(gnd), .vdd(vdd), .A(_20581_), .Y(_20581__bF_buf4) );
	BUFX4 BUFX4_1633 ( .gnd(gnd), .vdd(vdd), .A(_20581_), .Y(_20581__bF_buf3) );
	BUFX4 BUFX4_1634 ( .gnd(gnd), .vdd(vdd), .A(_20581_), .Y(_20581__bF_buf2) );
	BUFX4 BUFX4_1635 ( .gnd(gnd), .vdd(vdd), .A(_20581_), .Y(_20581__bF_buf1) );
	BUFX4 BUFX4_1636 ( .gnd(gnd), .vdd(vdd), .A(_20581_), .Y(_20581__bF_buf0) );
	BUFX4 BUFX4_1637 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf7) );
	BUFX4 BUFX4_1638 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf6) );
	BUFX4 BUFX4_1639 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf5) );
	BUFX4 BUFX4_1640 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf4) );
	BUFX4 BUFX4_1641 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf3) );
	BUFX4 BUFX4_1642 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf2) );
	BUFX4 BUFX4_1643 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf1) );
	BUFX4 BUFX4_1644 ( .gnd(gnd), .vdd(vdd), .A(_17371_), .Y(_17371__bF_buf0) );
	BUFX4 BUFX4_1645 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .Y(_4008__bF_buf5) );
	BUFX4 BUFX4_1646 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .Y(_4008__bF_buf4) );
	BUFX4 BUFX4_1647 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .Y(_4008__bF_buf3) );
	BUFX4 BUFX4_1648 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .Y(_4008__bF_buf2) );
	BUFX4 BUFX4_1649 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .Y(_4008__bF_buf1) );
	BUFX4 BUFX4_1650 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .Y(_4008__bF_buf0) );
	BUFX4 BUFX4_1651 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .Y(_5332__bF_buf3) );
	BUFX4 BUFX4_1652 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .Y(_5332__bF_buf2) );
	BUFX4 BUFX4_1653 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .Y(_5332__bF_buf1) );
	BUFX4 BUFX4_1654 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .Y(_5332__bF_buf0) );
	BUFX4 BUFX4_1655 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf10) );
	BUFX4 BUFX4_1656 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf9) );
	BUFX4 BUFX4_1657 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf8) );
	BUFX4 BUFX4_1658 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf7) );
	BUFX4 BUFX4_1659 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf6) );
	BUFX4 BUFX4_1660 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf5) );
	BUFX4 BUFX4_1661 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf4) );
	BUFX4 BUFX4_1662 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf3) );
	BUFX4 BUFX4_1663 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf2) );
	BUFX4 BUFX4_1664 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf1) );
	BUFX4 BUFX4_1665 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf0) );
	BUFX4 BUFX4_1666 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .Y(_3204__bF_buf4) );
	BUFX4 BUFX4_1667 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .Y(_3204__bF_buf3) );
	BUFX4 BUFX4_1668 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .Y(_3204__bF_buf2) );
	BUFX4 BUFX4_1669 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .Y(_3204__bF_buf1) );
	BUFX4 BUFX4_1670 ( .gnd(gnd), .vdd(vdd), .A(_3204_), .Y(_3204__bF_buf0) );
	BUFX4 BUFX4_1671 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf7) );
	BUFX4 BUFX4_1672 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf6) );
	BUFX4 BUFX4_1673 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf5) );
	BUFX4 BUFX4_1674 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf4) );
	BUFX4 BUFX4_1675 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf3) );
	BUFX4 BUFX4_1676 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf2) );
	BUFX4 BUFX4_1677 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf1) );
	BUFX4 BUFX4_1678 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .Y(_4100__bF_buf0) );
	BUFX4 BUFX4_1679 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf7) );
	BUFX4 BUFX4_1680 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf6) );
	BUFX4 BUFX4_1681 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf5) );
	BUFX4 BUFX4_1682 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf4) );
	BUFX4 BUFX4_1683 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf3) );
	BUFX4 BUFX4_1684 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf2) );
	BUFX4 BUFX4_1685 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf1) );
	BUFX4 BUFX4_1686 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .Y(_1768__bF_buf0) );
	BUFX4 BUFX4_1687 ( .gnd(gnd), .vdd(vdd), .A(_11776_), .Y(_11776__bF_buf3) );
	BUFX4 BUFX4_1688 ( .gnd(gnd), .vdd(vdd), .A(_11776_), .Y(_11776__bF_buf2) );
	BUFX4 BUFX4_1689 ( .gnd(gnd), .vdd(vdd), .A(_11776_), .Y(_11776__bF_buf1) );
	BUFX4 BUFX4_1690 ( .gnd(gnd), .vdd(vdd), .A(_11776_), .Y(_11776__bF_buf0) );
	BUFX4 BUFX4_1691 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_), .Y(aOperand_frameOut_17_bF_buf4) );
	BUFX4 BUFX4_1692 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_), .Y(aOperand_frameOut_17_bF_buf3) );
	BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_), .Y(aOperand_frameOut_17_bF_buf2) );
	BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_), .Y(aOperand_frameOut_17_bF_buf1) );
	BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_), .Y(aOperand_frameOut_17_bF_buf0) );
	BUFX4 BUFX4_1693 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .Y(_10676__bF_buf3) );
	BUFX4 BUFX4_1694 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .Y(_10676__bF_buf2) );
	BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .Y(_10676__bF_buf1) );
	BUFX4 BUFX4_1695 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .Y(_10676__bF_buf0) );
	BUFX4 BUFX4_1696 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf7) );
	BUFX4 BUFX4_1697 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf6) );
	BUFX4 BUFX4_1698 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf5) );
	BUFX4 BUFX4_1699 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf4) );
	BUFX4 BUFX4_1700 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf3) );
	BUFX4 BUFX4_1701 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf2) );
	BUFX4 BUFX4_1702 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf1) );
	BUFX4 BUFX4_1703 ( .gnd(gnd), .vdd(vdd), .A(_19432_), .Y(_19432__bF_buf0) );
	BUFX4 BUFX4_1704 ( .gnd(gnd), .vdd(vdd), .A(_17466_), .Y(_17466__bF_buf4) );
	BUFX4 BUFX4_1705 ( .gnd(gnd), .vdd(vdd), .A(_17466_), .Y(_17466__bF_buf3) );
	BUFX4 BUFX4_1706 ( .gnd(gnd), .vdd(vdd), .A(_17466_), .Y(_17466__bF_buf2) );
	BUFX4 BUFX4_1707 ( .gnd(gnd), .vdd(vdd), .A(_17466_), .Y(_17466__bF_buf1) );
	BUFX4 BUFX4_1708 ( .gnd(gnd), .vdd(vdd), .A(_17466_), .Y(_17466__bF_buf0) );
	BUFX4 BUFX4_1709 ( .gnd(gnd), .vdd(vdd), .A(_17436_), .Y(_17436__bF_buf4) );
	BUFX4 BUFX4_1710 ( .gnd(gnd), .vdd(vdd), .A(_17436_), .Y(_17436__bF_buf3) );
	BUFX4 BUFX4_1711 ( .gnd(gnd), .vdd(vdd), .A(_17436_), .Y(_17436__bF_buf2) );
	BUFX4 BUFX4_1712 ( .gnd(gnd), .vdd(vdd), .A(_17436_), .Y(_17436__bF_buf1) );
	BUFX4 BUFX4_1713 ( .gnd(gnd), .vdd(vdd), .A(_17436_), .Y(_17436__bF_buf0) );
	BUFX4 BUFX4_1714 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_), .Y(divider_absoluteValue_B_flipSign_result_22_bF_buf3) );
	BUFX4 BUFX4_1715 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_), .Y(divider_absoluteValue_B_flipSign_result_22_bF_buf2) );
	BUFX4 BUFX4_1716 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_), .Y(divider_absoluteValue_B_flipSign_result_22_bF_buf1) );
	BUFX4 BUFX4_1717 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_), .Y(divider_absoluteValue_B_flipSign_result_22_bF_buf0) );
	BUFX4 BUFX4_1718 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf7) );
	BUFX4 BUFX4_1719 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf6) );
	BUFX4 BUFX4_1720 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf5) );
	BUFX4 BUFX4_1721 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf4) );
	BUFX4 BUFX4_1722 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf3) );
	BUFX4 BUFX4_1723 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf2) );
	BUFX4 BUFX4_1724 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf1) );
	BUFX4 BUFX4_1725 ( .gnd(gnd), .vdd(vdd), .A(_20574_), .Y(_20574__bF_buf0) );
	BUFX4 BUFX4_1726 ( .gnd(gnd), .vdd(vdd), .A(_17394_), .Y(_17394__bF_buf4) );
	BUFX4 BUFX4_1727 ( .gnd(gnd), .vdd(vdd), .A(_17394_), .Y(_17394__bF_buf3) );
	BUFX4 BUFX4_1728 ( .gnd(gnd), .vdd(vdd), .A(_17394_), .Y(_17394__bF_buf2) );
	BUFX4 BUFX4_1729 ( .gnd(gnd), .vdd(vdd), .A(_17394_), .Y(_17394__bF_buf1) );
	BUFX4 BUFX4_1730 ( .gnd(gnd), .vdd(vdd), .A(_17394_), .Y(_17394__bF_buf0) );
	BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_), .Y(adder_bOperand_20_bF_buf3) );
	BUFX4 BUFX4_1731 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_), .Y(adder_bOperand_20_bF_buf2) );
	BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_), .Y(adder_bOperand_20_bF_buf1) );
	BUFX4 BUFX4_1732 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_), .Y(adder_bOperand_20_bF_buf0) );
	BUFX4 BUFX4_1733 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_), .Y(aOperand_frameOut_12_bF_buf4) );
	BUFX4 BUFX4_1734 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_), .Y(aOperand_frameOut_12_bF_buf3) );
	BUFX4 BUFX4_1735 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_), .Y(aOperand_frameOut_12_bF_buf2) );
	BUFX4 BUFX4_1736 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_), .Y(aOperand_frameOut_12_bF_buf1) );
	BUFX4 BUFX4_1737 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_), .Y(aOperand_frameOut_12_bF_buf0) );
	BUFX4 BUFX4_1738 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_), .Y(aOperand_frameOut_7_bF_buf4) );
	BUFX4 BUFX4_1739 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_), .Y(aOperand_frameOut_7_bF_buf3) );
	BUFX4 BUFX4_1740 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_), .Y(aOperand_frameOut_7_bF_buf2) );
	BUFX4 BUFX4_1741 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_), .Y(aOperand_frameOut_7_bF_buf1) );
	BUFX4 BUFX4_1742 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_), .Y(aOperand_frameOut_7_bF_buf0) );
	BUFX4 BUFX4_1743 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_), .Y(reg_dataIn_25_bF_buf4) );
	BUFX4 BUFX4_1744 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_), .Y(reg_dataIn_25_bF_buf3) );
	BUFX4 BUFX4_1745 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_), .Y(reg_dataIn_25_bF_buf2) );
	BUFX4 BUFX4_1746 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_), .Y(reg_dataIn_25_bF_buf1) );
	BUFX4 BUFX4_1747 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_), .Y(reg_dataIn_25_bF_buf0) );
	BUFX4 BUFX4_1748 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .Y(_5126__bF_buf3) );
	BUFX4 BUFX4_1749 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .Y(_5126__bF_buf2) );
	BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .Y(_5126__bF_buf1) );
	BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .Y(_5126__bF_buf0) );
	BUFX4 BUFX4_1750 ( .gnd(gnd), .vdd(vdd), .A(_20611_), .Y(_20611__bF_buf4) );
	BUFX4 BUFX4_1751 ( .gnd(gnd), .vdd(vdd), .A(_20611_), .Y(_20611__bF_buf3) );
	BUFX4 BUFX4_1752 ( .gnd(gnd), .vdd(vdd), .A(_20611_), .Y(_20611__bF_buf2) );
	BUFX4 BUFX4_1753 ( .gnd(gnd), .vdd(vdd), .A(_20611_), .Y(_20611__bF_buf1) );
	BUFX4 BUFX4_1754 ( .gnd(gnd), .vdd(vdd), .A(_20611_), .Y(_20611__bF_buf0) );
	BUFX4 BUFX4_1755 ( .gnd(gnd), .vdd(vdd), .A(_17461_), .Y(_17461__bF_buf4) );
	BUFX4 BUFX4_1756 ( .gnd(gnd), .vdd(vdd), .A(_17461_), .Y(_17461__bF_buf3) );
	BUFX4 BUFX4_1757 ( .gnd(gnd), .vdd(vdd), .A(_17461_), .Y(_17461__bF_buf2) );
	BUFX4 BUFX4_1758 ( .gnd(gnd), .vdd(vdd), .A(_17461_), .Y(_17461__bF_buf1) );
	BUFX4 BUFX4_1759 ( .gnd(gnd), .vdd(vdd), .A(_17461_), .Y(_17461__bF_buf0) );
	BUFX4 BUFX4_1760 ( .gnd(gnd), .vdd(vdd), .A(_17431_), .Y(_17431__bF_buf4) );
	BUFX4 BUFX4_1761 ( .gnd(gnd), .vdd(vdd), .A(_17431_), .Y(_17431__bF_buf3) );
	BUFX4 BUFX4_1762 ( .gnd(gnd), .vdd(vdd), .A(_17431_), .Y(_17431__bF_buf2) );
	BUFX4 BUFX4_1763 ( .gnd(gnd), .vdd(vdd), .A(_17431_), .Y(_17431__bF_buf1) );
	BUFX4 BUFX4_1764 ( .gnd(gnd), .vdd(vdd), .A(_17431_), .Y(_17431__bF_buf0) );
	BUFX4 BUFX4_1765 ( .gnd(gnd), .vdd(vdd), .A(_17401_), .Y(_17401__bF_buf4) );
	BUFX4 BUFX4_1766 ( .gnd(gnd), .vdd(vdd), .A(_17401_), .Y(_17401__bF_buf3) );
	BUFX4 BUFX4_1767 ( .gnd(gnd), .vdd(vdd), .A(_17401_), .Y(_17401__bF_buf2) );
	BUFX4 BUFX4_1768 ( .gnd(gnd), .vdd(vdd), .A(_17401_), .Y(_17401__bF_buf1) );
	BUFX4 BUFX4_1769 ( .gnd(gnd), .vdd(vdd), .A(_17401_), .Y(_17401__bF_buf0) );
	BUFX4 BUFX4_1770 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip), .Y(divider_absoluteValue_B_flipSign_flip_bF_buf5) );
	BUFX4 BUFX4_1771 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip), .Y(divider_absoluteValue_B_flipSign_flip_bF_buf4) );
	BUFX4 BUFX4_1772 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip), .Y(divider_absoluteValue_B_flipSign_flip_bF_buf3) );
	BUFX4 BUFX4_1773 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip), .Y(divider_absoluteValue_B_flipSign_flip_bF_buf2) );
	BUFX4 BUFX4_1774 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip), .Y(divider_absoluteValue_B_flipSign_flip_bF_buf1) );
	BUFX4 BUFX4_1775 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip), .Y(divider_absoluteValue_B_flipSign_flip_bF_buf0) );
	BUFX4 BUFX4_1776 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_), .Y(aOperand_frameOut_2_bF_buf4) );
	BUFX4 BUFX4_1777 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_), .Y(aOperand_frameOut_2_bF_buf3) );
	BUFX4 BUFX4_1778 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_), .Y(aOperand_frameOut_2_bF_buf2) );
	BUFX4 BUFX4_1779 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_), .Y(aOperand_frameOut_2_bF_buf1) );
	BUFX4 BUFX4_1780 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_), .Y(aOperand_frameOut_2_bF_buf0) );
	BUFX4 BUFX4_1781 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_), .Y(reg_dataIn_20_bF_buf4) );
	BUFX4 BUFX4_1782 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_), .Y(reg_dataIn_20_bF_buf3) );
	BUFX4 BUFX4_1783 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_), .Y(reg_dataIn_20_bF_buf2) );
	BUFX4 BUFX4_1784 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_), .Y(reg_dataIn_20_bF_buf1) );
	BUFX4 BUFX4_1785 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_), .Y(reg_dataIn_20_bF_buf0) );
	BUFX4 BUFX4_1786 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .Y(_2229__bF_buf4) );
	BUFX4 BUFX4_1787 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .Y(_2229__bF_buf3) );
	BUFX4 BUFX4_1788 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .Y(_2229__bF_buf2) );
	BUFX4 BUFX4_1789 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .Y(_2229__bF_buf1) );
	BUFX4 BUFX4_1790 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .Y(_2229__bF_buf0) );
	BUFX4 BUFX4_1791 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .Y(_4424__bF_buf3) );
	BUFX4 BUFX4_1792 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .Y(_4424__bF_buf2) );
	BUFX4 BUFX4_1793 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .Y(_4424__bF_buf1) );
	BUFX4 BUFX4_1794 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .Y(_4424__bF_buf0) );
	BUFX4 BUFX4_1795 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf7) );
	BUFX4 BUFX4_1796 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf6) );
	BUFX4 BUFX4_1797 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf5) );
	BUFX4 BUFX4_1798 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf4) );
	BUFX4 BUFX4_1799 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf3) );
	BUFX4 BUFX4_1800 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf2) );
	BUFX4 BUFX4_1801 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf1) );
	BUFX4 BUFX4_1802 ( .gnd(gnd), .vdd(vdd), .A(_19328_), .Y(_19328__bF_buf0) );
	BUFX4 BUFX4_1803 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_), .Y(adder_bOperand_18_bF_buf3) );
	BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_), .Y(adder_bOperand_18_bF_buf2) );
	BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_), .Y(adder_bOperand_18_bF_buf1) );
	BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_), .Y(adder_bOperand_18_bF_buf0) );
	BUFX4 BUFX4_1804 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf7) );
	BUFX4 BUFX4_1805 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf6) );
	BUFX4 BUFX4_1806 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf5) );
	BUFX4 BUFX4_1807 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf4) );
	BUFX4 BUFX4_1808 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf3) );
	BUFX4 BUFX4_1809 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf2) );
	BUFX4 BUFX4_1810 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf1) );
	BUFX4 BUFX4_1811 ( .gnd(gnd), .vdd(vdd), .A(_19256_), .Y(_19256__bF_buf0) );
	BUFX4 BUFX4_1812 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_), .Y(reg_dataIn_8_bF_buf4) );
	BUFX4 BUFX4_1813 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_), .Y(reg_dataIn_8_bF_buf3) );
	BUFX4 BUFX4_1814 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_), .Y(reg_dataIn_8_bF_buf2) );
	BUFX4 BUFX4_1815 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_), .Y(reg_dataIn_8_bF_buf1) );
	BUFX4 BUFX4_1816 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_), .Y(reg_dataIn_8_bF_buf0) );
	BUFX4 BUFX4_1817 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf7) );
	BUFX4 BUFX4_1818 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf6) );
	BUFX4 BUFX4_1819 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf5) );
	BUFX4 BUFX4_1820 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf4) );
	BUFX4 BUFX4_1821 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf3) );
	BUFX4 BUFX4_1822 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf2) );
	BUFX4 BUFX4_1823 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf1) );
	BUFX4 BUFX4_1824 ( .gnd(gnd), .vdd(vdd), .A(_20296_), .Y(_20296__bF_buf0) );
	BUFX4 BUFX4_1825 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_), .Y(divider_absoluteValue_B_flipSign_result_15_bF_buf4) );
	BUFX4 BUFX4_1826 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_), .Y(divider_absoluteValue_B_flipSign_result_15_bF_buf3) );
	BUFX4 BUFX4_1827 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_), .Y(divider_absoluteValue_B_flipSign_result_15_bF_buf2) );
	BUFX4 BUFX4_1828 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_), .Y(divider_absoluteValue_B_flipSign_result_15_bF_buf1) );
	BUFX4 BUFX4_1829 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_), .Y(divider_absoluteValue_B_flipSign_result_15_bF_buf0) );
	BUFX4 BUFX4_1830 ( .gnd(gnd), .vdd(vdd), .A(_20567_), .Y(_20567__bF_buf4) );
	BUFX4 BUFX4_1831 ( .gnd(gnd), .vdd(vdd), .A(_20567_), .Y(_20567__bF_buf3) );
	BUFX4 BUFX4_1832 ( .gnd(gnd), .vdd(vdd), .A(_20567_), .Y(_20567__bF_buf2) );
	BUFX4 BUFX4_1833 ( .gnd(gnd), .vdd(vdd), .A(_20567_), .Y(_20567__bF_buf1) );
	BUFX4 BUFX4_1834 ( .gnd(gnd), .vdd(vdd), .A(_20567_), .Y(_20567__bF_buf0) );
	BUFX4 BUFX4_1835 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_), .Y(adder_bOperand_13_bF_buf3) );
	BUFX4 BUFX4_1836 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_), .Y(adder_bOperand_13_bF_buf2) );
	BUFX4 BUFX4_1837 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_), .Y(adder_bOperand_13_bF_buf1) );
	BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_), .Y(adder_bOperand_13_bF_buf0) );
	BUFX4 BUFX4_1838 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_), .Y(reg_dataIn_3_bF_buf4) );
	BUFX4 BUFX4_1839 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_), .Y(reg_dataIn_3_bF_buf3) );
	BUFX4 BUFX4_1840 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_), .Y(reg_dataIn_3_bF_buf2) );
	BUFX4 BUFX4_1841 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_), .Y(reg_dataIn_3_bF_buf1) );
	BUFX4 BUFX4_1842 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_), .Y(reg_dataIn_3_bF_buf0) );
	BUFX4 BUFX4_1843 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_), .Y(reg_dataIn_18_bF_buf4) );
	BUFX4 BUFX4_1844 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_), .Y(reg_dataIn_18_bF_buf3) );
	BUFX4 BUFX4_1845 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_), .Y(reg_dataIn_18_bF_buf2) );
	BUFX4 BUFX4_1846 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_), .Y(reg_dataIn_18_bF_buf1) );
	BUFX4 BUFX4_1847 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_), .Y(reg_dataIn_18_bF_buf0) );
	BUFX4 BUFX4_1848 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf4) );
	BUFX4 BUFX4_1849 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf3) );
	BUFX4 BUFX4_1850 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf2) );
	BUFX4 BUFX4_1851 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf1) );
	BUFX4 BUFX4_1852 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .Y(_11560__bF_buf0) );
	BUFX4 BUFX4_1853 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf6) );
	BUFX4 BUFX4_1854 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf5) );
	BUFX4 BUFX4_1855 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf4) );
	BUFX4 BUFX4_1856 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf3) );
	BUFX4 BUFX4_1857 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf2) );
	BUFX4 BUFX4_1858 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf1) );
	BUFX4 BUFX4_1859 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_), .Y(divider_absoluteValue_B_flipSign_result_8_bF_buf0) );
	BUFX4 BUFX4_1860 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf7) );
	BUFX4 BUFX4_1861 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf6) );
	BUFX4 BUFX4_1862 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf5) );
	BUFX4 BUFX4_1863 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf4) );
	BUFX4 BUFX4_1864 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf3) );
	BUFX4 BUFX4_1865 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf2) );
	BUFX4 BUFX4_1866 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf1) );
	BUFX4 BUFX4_1867 ( .gnd(gnd), .vdd(vdd), .A(_20002_), .Y(_20002__bF_buf0) );
	BUFX4 BUFX4_1868 ( .gnd(gnd), .vdd(vdd), .A(_17454_), .Y(_17454__bF_buf4) );
	BUFX4 BUFX4_1869 ( .gnd(gnd), .vdd(vdd), .A(_17454_), .Y(_17454__bF_buf3) );
	BUFX4 BUFX4_1870 ( .gnd(gnd), .vdd(vdd), .A(_17454_), .Y(_17454__bF_buf2) );
	BUFX4 BUFX4_1871 ( .gnd(gnd), .vdd(vdd), .A(_17454_), .Y(_17454__bF_buf1) );
	BUFX4 BUFX4_1872 ( .gnd(gnd), .vdd(vdd), .A(_17454_), .Y(_17454__bF_buf0) );
	BUFX4 BUFX4_1873 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_), .Y(divider_absoluteValue_B_flipSign_result_10_bF_buf5) );
	BUFX4 BUFX4_1874 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_), .Y(divider_absoluteValue_B_flipSign_result_10_bF_buf4) );
	BUFX4 BUFX4_1875 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_), .Y(divider_absoluteValue_B_flipSign_result_10_bF_buf3) );
	BUFX4 BUFX4_1876 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_), .Y(divider_absoluteValue_B_flipSign_result_10_bF_buf2) );
	BUFX4 BUFX4_1877 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_), .Y(divider_absoluteValue_B_flipSign_result_10_bF_buf1) );
	BUFX4 BUFX4_1878 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_), .Y(divider_absoluteValue_B_flipSign_result_10_bF_buf0) );
	BUFX4 BUFX4_1879 ( .gnd(gnd), .vdd(vdd), .A(_20562_), .Y(_20562__bF_buf5) );
	BUFX4 BUFX4_1880 ( .gnd(gnd), .vdd(vdd), .A(_20562_), .Y(_20562__bF_buf4) );
	BUFX4 BUFX4_1881 ( .gnd(gnd), .vdd(vdd), .A(_20562_), .Y(_20562__bF_buf3) );
	BUFX4 BUFX4_1882 ( .gnd(gnd), .vdd(vdd), .A(_20562_), .Y(_20562__bF_buf2) );
	BUFX4 BUFX4_1883 ( .gnd(gnd), .vdd(vdd), .A(_20562_), .Y(_20562__bF_buf1) );
	BUFX4 BUFX4_1884 ( .gnd(gnd), .vdd(vdd), .A(_20562_), .Y(_20562__bF_buf0) );
	BUFX4 BUFX4_1885 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_), .Y(adder_bOperand_9_bF_buf4) );
	BUFX4 BUFX4_1886 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_), .Y(adder_bOperand_9_bF_buf3) );
	BUFX4 BUFX4_1887 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_), .Y(adder_bOperand_9_bF_buf2) );
	BUFX4 BUFX4_1888 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_), .Y(adder_bOperand_9_bF_buf1) );
	BUFX4 BUFX4_1889 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_), .Y(adder_bOperand_9_bF_buf0) );
	BUFX4 BUFX4_1890 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf7) );
	BUFX4 BUFX4_1891 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf6) );
	BUFX4 BUFX4_1892 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf5) );
	BUFX4 BUFX4_1893 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf4) );
	BUFX4 BUFX4_1894 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf3) );
	BUFX4 BUFX4_1895 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf2) );
	BUFX4 BUFX4_1896 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf1) );
	BUFX4 BUFX4_1897 ( .gnd(gnd), .vdd(vdd), .A(_20231_), .Y(_20231__bF_buf0) );
	BUFX4 BUFX4_1898 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip), .Y(divider_divFlip_bF_buf5) );
	BUFX4 BUFX4_1899 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip), .Y(divider_divFlip_bF_buf4) );
	BUFX4 BUFX4_1900 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip), .Y(divider_divFlip_bF_buf3) );
	BUFX4 BUFX4_1901 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip), .Y(divider_divFlip_bF_buf2) );
	BUFX4 BUFX4_1902 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip), .Y(divider_divFlip_bF_buf1) );
	BUFX4 BUFX4_1903 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip), .Y(divider_divFlip_bF_buf0) );
	BUFX4 BUFX4_1904 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_), .Y(reg_dataIn_13_bF_buf4) );
	BUFX4 BUFX4_1905 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_), .Y(reg_dataIn_13_bF_buf3) );
	BUFX4 BUFX4_1906 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_), .Y(reg_dataIn_13_bF_buf2) );
	BUFX4 BUFX4_1907 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_), .Y(reg_dataIn_13_bF_buf1) );
	BUFX4 BUFX4_1908 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_), .Y(reg_dataIn_13_bF_buf0) );
	BUFX4 BUFX4_1909 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_), .Y(divider_divuResult_16_bF_buf5) );
	BUFX4 BUFX4_1910 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_), .Y(divider_divuResult_16_bF_buf4) );
	BUFX4 BUFX4_1911 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_), .Y(divider_divuResult_16_bF_buf3) );
	BUFX4 BUFX4_1912 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_), .Y(divider_divuResult_16_bF_buf2) );
	BUFX4 BUFX4_1913 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_), .Y(divider_divuResult_16_bF_buf1) );
	BUFX4 BUFX4_1914 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_), .Y(divider_divuResult_16_bF_buf0) );
	BUFX4 BUFX4_1915 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf7) );
	BUFX4 BUFX4_1916 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf6) );
	BUFX4 BUFX4_1917 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf5) );
	BUFX4 BUFX4_1918 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf4) );
	BUFX4 BUFX4_1919 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf3) );
	BUFX4 BUFX4_1920 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf2) );
	BUFX4 BUFX4_1921 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf1) );
	BUFX4 BUFX4_1922 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_), .Y(divider_absoluteValue_B_flipSign_result_3_bF_buf0) );
	BUFX4 BUFX4_1923 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_), .Y(adder_bOperand_4_bF_buf5) );
	BUFX4 BUFX4_1924 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_), .Y(adder_bOperand_4_bF_buf4) );
	BUFX4 BUFX4_1925 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_), .Y(adder_bOperand_4_bF_buf3) );
	BUFX4 BUFX4_1926 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_), .Y(adder_bOperand_4_bF_buf2) );
	BUFX4 BUFX4_1927 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_), .Y(adder_bOperand_4_bF_buf1) );
	BUFX4 BUFX4_1928 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_), .Y(adder_bOperand_4_bF_buf0) );
	BUFX4 BUFX4_1929 ( .gnd(gnd), .vdd(vdd), .A(_14684_), .Y(_14684__bF_buf3) );
	BUFX4 BUFX4_1930 ( .gnd(gnd), .vdd(vdd), .A(_14684_), .Y(_14684__bF_buf2) );
	BUFX4 BUFX4_1931 ( .gnd(gnd), .vdd(vdd), .A(_14684_), .Y(_14684__bF_buf1) );
	BUFX4 BUFX4_1932 ( .gnd(gnd), .vdd(vdd), .A(_14684_), .Y(_14684__bF_buf0) );
	BUFX4 BUFX4_1933 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_), .Y(divider_divuResult_11_bF_buf5) );
	BUFX4 BUFX4_1934 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_), .Y(divider_divuResult_11_bF_buf4) );
	BUFX4 BUFX4_1935 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_), .Y(divider_divuResult_11_bF_buf3) );
	BUFX4 BUFX4_1936 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_), .Y(divider_divuResult_11_bF_buf2) );
	BUFX4 BUFX4_1937 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_), .Y(divider_divuResult_11_bF_buf1) );
	BUFX4 BUFX4_1938 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_), .Y(divider_divuResult_11_bF_buf0) );
	BUFX4 BUFX4_1939 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf6) );
	BUFX4 BUFX4_1940 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf5) );
	BUFX4 BUFX4_1941 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf4) );
	BUFX4 BUFX4_1942 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf3) );
	BUFX4 BUFX4_1943 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf2) );
	BUFX4 BUFX4_1944 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf1) );
	BUFX4 BUFX4_1945 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_), .Y(divider_divuResult_7_bF_buf0) );
	BUFX4 BUFX4_1946 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf7) );
	BUFX4 BUFX4_1947 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf6) );
	BUFX4 BUFX4_1948 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf5) );
	BUFX4 BUFX4_1949 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf4) );
	BUFX4 BUFX4_1950 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf3) );
	BUFX4 BUFX4_1951 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf2) );
	BUFX4 BUFX4_1952 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf1) );
	BUFX4 BUFX4_1953 ( .gnd(gnd), .vdd(vdd), .A(_20458_), .Y(_20458__bF_buf0) );
	BUFX4 BUFX4_1954 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf6) );
	BUFX4 BUFX4_1955 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf5) );
	BUFX4 BUFX4_1956 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf4) );
	BUFX4 BUFX4_1957 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf3) );
	BUFX4 BUFX4_1958 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf2) );
	BUFX4 BUFX4_1959 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf1) );
	BUFX4 BUFX4_1960 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_), .Y(bLoc_frameOut_4_bF_buf0) );
	BUFX4 BUFX4_1961 ( .gnd(gnd), .vdd(vdd), .A(_11252_), .Y(_11252__bF_buf4) );
	BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(_11252_), .Y(_11252__bF_buf3) );
	BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(_11252_), .Y(_11252__bF_buf2) );
	BUFX4 BUFX4_1962 ( .gnd(gnd), .vdd(vdd), .A(_11252_), .Y(_11252__bF_buf1) );
	BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(_11252_), .Y(_11252__bF_buf0) );
	BUFX4 BUFX4_1963 ( .gnd(gnd), .vdd(vdd), .A(_20585_), .Y(_20585__bF_buf4) );
	BUFX4 BUFX4_1964 ( .gnd(gnd), .vdd(vdd), .A(_20585_), .Y(_20585__bF_buf3) );
	BUFX4 BUFX4_1965 ( .gnd(gnd), .vdd(vdd), .A(_20585_), .Y(_20585__bF_buf2) );
	BUFX4 BUFX4_1966 ( .gnd(gnd), .vdd(vdd), .A(_20585_), .Y(_20585__bF_buf1) );
	BUFX4 BUFX4_1967 ( .gnd(gnd), .vdd(vdd), .A(_20585_), .Y(_20585__bF_buf0) );
	BUFX4 BUFX4_1968 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf7) );
	BUFX4 BUFX4_1969 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf6) );
	BUFX4 BUFX4_1970 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf5) );
	BUFX4 BUFX4_1971 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf4) );
	BUFX4 BUFX4_1972 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf3) );
	BUFX4 BUFX4_1973 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf2) );
	BUFX4 BUFX4_1974 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf1) );
	BUFX4 BUFX4_1975 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_), .Y(divider_divuResult_2_bF_buf0) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeEnable_out), .B(frameWriteController_result_we), .Y(registers_writeEnable) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_0_), .Y(_0_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_0_), .B(immediateSelect_frameOut_bF_buf7), .Y(_1_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_0_), .C(_1_), .Y(bOperand_frameIn_0_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_1_), .Y(_2_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_1_), .Y(_3_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_2_), .C(_3_), .Y(bOperand_frameIn_1_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_2_), .Y(_4_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_2_), .Y(_5_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_4_), .C(_5_), .Y(bOperand_frameIn_2_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_3_), .Y(_6_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_3_), .Y(_7_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_6_), .C(_7_), .Y(bOperand_frameIn_3_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_4_), .Y(_8_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_4_), .Y(_9_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_8_), .C(_9_), .Y(bOperand_frameIn_4_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_5_), .Y(_10_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_5_), .Y(_11_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_10_), .C(_11_), .Y(bOperand_frameIn_5_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_6_), .Y(_12_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_6_), .Y(_13_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_12_), .C(_13_), .Y(bOperand_frameIn_6_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_7_), .Y(_14_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_7_), .Y(_15_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_14_), .C(_15_), .Y(bOperand_frameIn_7_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_8_), .Y(_16_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_8_), .Y(_17_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_16_), .C(_17_), .Y(bOperand_frameIn_8_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_9_), .Y(_18_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_9_), .Y(_19_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_18_), .C(_19_), .Y(bOperand_frameIn_9_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_10_), .Y(_20_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_10_), .Y(_21_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_20_), .C(_21_), .Y(bOperand_frameIn_10_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_11_), .Y(_22_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_11_), .Y(_23_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_22_), .C(_23_), .Y(bOperand_frameIn_11_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_12_), .Y(_24_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_12_), .Y(_25_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_24_), .C(_25_), .Y(bOperand_frameIn_12_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_13_), .Y(_26_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_13_), .Y(_27_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_26_), .C(_27_), .Y(bOperand_frameIn_13_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_14_), .Y(_28_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_14_), .Y(_29_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_28_), .C(_29_), .Y(bOperand_frameIn_14_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_15_), .Y(_30_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_15_), .Y(_31_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_30_), .C(_31_), .Y(bOperand_frameIn_15_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_16_), .Y(_32_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_16_), .Y(_33_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_32_), .C(_33_), .Y(bOperand_frameIn_16_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_17_), .Y(_34_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_17_), .Y(_35_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_34_), .C(_35_), .Y(bOperand_frameIn_17_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_18_), .Y(_36_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_18_), .Y(_37_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_36_), .C(_37_), .Y(bOperand_frameIn_18_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_19_), .Y(_38_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_19_), .Y(_39_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_38_), .C(_39_), .Y(bOperand_frameIn_19_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_20_), .Y(_40_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_20_), .Y(_41_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_40_), .C(_41_), .Y(bOperand_frameIn_20_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_21_), .Y(_42_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_21_), .Y(_43_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_42_), .C(_43_), .Y(bOperand_frameIn_21_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_22_), .Y(_44_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_22_), .Y(_45_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_44_), .C(_45_), .Y(bOperand_frameIn_22_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_23_), .Y(_46_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_23_), .Y(_47_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_46_), .C(_47_), .Y(bOperand_frameIn_23_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_24_), .Y(_48_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_24_), .Y(_49_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_48_), .C(_49_), .Y(bOperand_frameIn_24_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_25_), .Y(_50_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_25_), .Y(_51_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_50_), .C(_51_), .Y(bOperand_frameIn_25_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_26_), .Y(_52_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_26_), .Y(_53_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_52_), .C(_53_), .Y(bOperand_frameIn_26_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_27_), .Y(_54_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_27_), .Y(_55_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_54_), .C(_55_), .Y(bOperand_frameIn_27_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_28_), .Y(_56_) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(immediateVal_frameOut_28_), .Y(_57_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf6), .B(_56_), .C(_57_), .Y(bOperand_frameIn_28_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_29_), .Y(_58_) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf5), .B(immediateVal_frameOut_29_), .Y(_59_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf4), .B(_58_), .C(_59_), .Y(bOperand_frameIn_29_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_30_), .Y(_60_) );
	NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf3), .B(immediateVal_frameOut_30_), .Y(_61_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf2), .B(_60_), .C(_61_), .Y(bOperand_frameIn_30_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(readB_regOut_31_), .Y(_62_) );
	NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf1), .B(immediateVal_frameOut_31_), .Y(_63_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf0), .B(_62_), .C(_63_), .Y(bOperand_frameIn_31_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_1_), .Y(_64_) );
	NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_0_), .B(_64_), .Y(_65_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_2_), .B(_65_), .Y(_66_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(comparator_equal_0_), .Y(_67_) );
	INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_2_), .Y(_68_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_1_), .B(instructionFrame_resultSelect_out_0_), .Y(_69_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_0_), .C(_69__bF_buf4), .Y(_70_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_2_), .B(instructionFrame_resultSelect_out_0_), .C(_64_), .Y(_71_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_71__bF_buf4), .C(_70_), .Y(_72_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(mulOut_0_), .B(_66__bF_buf4), .C(_72_), .Y(_73_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_0_), .Y(_74_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(comparator_greater_0_), .Y(_75_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_0_), .Y(_76_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_2_), .B(_64_), .C(_76_), .Y(_77_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_1_), .B(instructionFrame_resultSelect_out_0_), .C(_68__bF_buf3), .Y(_78_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_78__bF_buf4), .C(_75_), .D(_77__bF_buf4), .Y(_79_) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(comparator_less_0_), .Y(_80_) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(divideOut_0_), .Y(_81_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_1_), .B(_68__bF_buf2), .C(_76_), .Y(_82_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_2_), .B(instructionFrame_resultSelect_out_1_), .C(_76_), .Y(_83_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_83__bF_buf4), .C(_81_), .D(_82__bF_buf4), .Y(_84_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_84_), .Y(_85_) );
	NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_85_), .Y(reg_dataIn_0_) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_86_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_1_), .C(_69__bF_buf3), .Y(_87_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_71__bF_buf3), .C(_87_), .Y(_88_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(mulOut_1_), .B(_66__bF_buf3), .C(_88_), .Y(_89_) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_1_), .Y(_90_) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_91_) );
	OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_78__bF_buf3), .C(_91_), .D(_77__bF_buf3), .Y(_92_) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_93_) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(divideOut_1_), .Y(_94_) );
	OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_83__bF_buf3), .C(_94_), .D(_82__bF_buf3), .Y(_95_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_95_), .Y(_96_) );
	NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_96_), .Y(reg_dataIn_1_) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_97_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(adder_result_2_), .C(_69__bF_buf2), .Y(_98_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_71__bF_buf2), .C(_98_), .Y(_99_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(mulOut_2_), .B(_66__bF_buf2), .C(_99_), .Y(_100_) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_2_), .Y(_101_) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_102_) );
	OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_78__bF_buf2), .C(_102_), .D(_77__bF_buf2), .Y(_103_) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_104_) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(divideOut_2_), .Y(_105_) );
	OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_83__bF_buf2), .C(_105_), .D(_82__bF_buf2), .Y(_106_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_106_), .Y(_107_) );
	NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_107_), .Y(reg_dataIn_2_) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_108_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_3_), .C(_69__bF_buf1), .Y(_109_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_71__bF_buf1), .C(_109_), .Y(_110_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(mulOut_3_), .B(_66__bF_buf1), .C(_110_), .Y(_111_) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_3_), .Y(_112_) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_113_) );
	OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_78__bF_buf1), .C(_113_), .D(_77__bF_buf1), .Y(_114_) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_115_) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(divideOut_3_), .Y(_116_) );
	OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_83__bF_buf1), .C(_116_), .D(_82__bF_buf1), .Y(_117_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_117_), .Y(_118_) );
	NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_118_), .Y(reg_dataIn_3_) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_119_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(adder_result_4_), .C(_69__bF_buf0), .Y(_120_) );
	OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_71__bF_buf0), .C(_120_), .Y(_121_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(mulOut_4_), .B(_66__bF_buf0), .C(_121_), .Y(_122_) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_4_), .Y(_123_) );
	INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_124_) );
	OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_78__bF_buf0), .C(_124_), .D(_77__bF_buf0), .Y(_125_) );
	INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_126_) );
	INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(divideOut_4_), .Y(_127_) );
	OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_83__bF_buf0), .C(_127_), .D(_82__bF_buf0), .Y(_128_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_128_), .Y(_129_) );
	NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_129_), .Y(reg_dataIn_4_) );
	INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_130_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(adder_result_5_), .C(_69__bF_buf4), .Y(_131_) );
	OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_71__bF_buf4), .C(_131_), .Y(_132_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(mulOut_5_), .B(_66__bF_buf4), .C(_132_), .Y(_133_) );
	INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_5_), .Y(_134_) );
	INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_135_) );
	OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_78__bF_buf4), .C(_135_), .D(_77__bF_buf4), .Y(_136_) );
	INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_137_) );
	INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(divideOut_5_), .Y(_138_) );
	OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_83__bF_buf4), .C(_138_), .D(_82__bF_buf4), .Y(_139_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_139_), .Y(_140_) );
	NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_140_), .Y(reg_dataIn_5_) );
	INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_141_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_6_), .C(_69__bF_buf3), .Y(_142_) );
	OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_71__bF_buf3), .C(_142_), .Y(_143_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(mulOut_6_), .B(_66__bF_buf3), .C(_143_), .Y(_144_) );
	INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_6_), .Y(_145_) );
	INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_146_) );
	OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_78__bF_buf3), .C(_146_), .D(_77__bF_buf3), .Y(_147_) );
	INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_148_) );
	INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(divideOut_6_), .Y(_149_) );
	OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_83__bF_buf3), .C(_149_), .D(_82__bF_buf3), .Y(_150_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_150_), .Y(_151_) );
	NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_151_), .Y(reg_dataIn_6_) );
	INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_152_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(adder_result_7_), .C(_69__bF_buf2), .Y(_153_) );
	OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_71__bF_buf2), .C(_153_), .Y(_154_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(mulOut_7_), .B(_66__bF_buf2), .C(_154_), .Y(_155_) );
	INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_7_), .Y(_156_) );
	INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_157_) );
	OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_78__bF_buf2), .C(_157_), .D(_77__bF_buf2), .Y(_158_) );
	INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_159_) );
	INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(divideOut_7_), .Y(_160_) );
	OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_83__bF_buf2), .C(_160_), .D(_82__bF_buf2), .Y(_161_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_161_), .Y(_162_) );
	NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_162_), .Y(reg_dataIn_7_) );
	INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_163_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_8_), .C(_69__bF_buf1), .Y(_164_) );
	OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_71__bF_buf1), .C(_164_), .Y(_165_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(mulOut_8_), .B(_66__bF_buf1), .C(_165_), .Y(_166_) );
	INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_8_), .Y(_167_) );
	INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_168_) );
	OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_78__bF_buf1), .C(_168_), .D(_77__bF_buf1), .Y(_169_) );
	INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_170_) );
	INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(divideOut_8_), .Y(_171_) );
	OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_83__bF_buf1), .C(_171_), .D(_82__bF_buf1), .Y(_172_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_172_), .Y(_173_) );
	NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_173_), .Y(reg_dataIn_8_) );
	INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_174_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(adder_result_9_), .C(_69__bF_buf0), .Y(_175_) );
	OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_71__bF_buf0), .C(_175_), .Y(_176_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(mulOut_9_), .B(_66__bF_buf0), .C(_176_), .Y(_177_) );
	INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_9_), .Y(_178_) );
	INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_179_) );
	OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_78__bF_buf0), .C(_179_), .D(_77__bF_buf0), .Y(_180_) );
	INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_181_) );
	INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(divideOut_9_), .Y(_182_) );
	OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_83__bF_buf0), .C(_182_), .D(_82__bF_buf0), .Y(_183_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_183_), .Y(_184_) );
	NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_184_), .Y(reg_dataIn_9_) );
	INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_185_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(adder_result_10_), .C(_69__bF_buf4), .Y(_186_) );
	OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_71__bF_buf4), .C(_186_), .Y(_187_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(mulOut_10_), .B(_66__bF_buf4), .C(_187_), .Y(_188_) );
	INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_10_), .Y(_189_) );
	INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_190_) );
	OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_78__bF_buf4), .C(_190_), .D(_77__bF_buf4), .Y(_191_) );
	INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_192_) );
	INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(divideOut_10_), .Y(_193_) );
	OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_83__bF_buf4), .C(_193_), .D(_82__bF_buf4), .Y(_194_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_194_), .Y(_195_) );
	NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_195_), .Y(reg_dataIn_10_) );
	INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_196_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_11_), .C(_69__bF_buf3), .Y(_197_) );
	OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_71__bF_buf3), .C(_197_), .Y(_198_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(mulOut_11_), .B(_66__bF_buf3), .C(_198_), .Y(_199_) );
	INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_11_), .Y(_200_) );
	INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_201_) );
	OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_78__bF_buf3), .C(_201_), .D(_77__bF_buf3), .Y(_202_) );
	INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_203_) );
	INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(divideOut_11_), .Y(_204_) );
	OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_83__bF_buf3), .C(_204_), .D(_82__bF_buf3), .Y(_205_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_205_), .Y(_206_) );
	NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_206_), .Y(reg_dataIn_11_) );
	INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_207_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(adder_result_12_), .C(_69__bF_buf2), .Y(_208_) );
	OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_71__bF_buf2), .C(_208_), .Y(_209_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(mulOut_12_), .B(_66__bF_buf2), .C(_209_), .Y(_210_) );
	INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_12_), .Y(_211_) );
	INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_212_) );
	OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_78__bF_buf2), .C(_212_), .D(_77__bF_buf2), .Y(_213_) );
	INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_214_) );
	INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(divideOut_12_), .Y(_215_) );
	OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_83__bF_buf2), .C(_215_), .D(_82__bF_buf2), .Y(_216_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_216_), .Y(_217_) );
	NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_217_), .Y(reg_dataIn_12_) );
	INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_218_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_13_), .C(_69__bF_buf1), .Y(_219_) );
	OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_71__bF_buf1), .C(_219_), .Y(_220_) );
	AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(mulOut_13_), .B(_66__bF_buf1), .C(_220_), .Y(_221_) );
	INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_13_), .Y(_222_) );
	INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_223_) );
	OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_78__bF_buf1), .C(_223_), .D(_77__bF_buf1), .Y(_224_) );
	INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_225_) );
	INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(divideOut_13_), .Y(_226_) );
	OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_83__bF_buf1), .C(_226_), .D(_82__bF_buf1), .Y(_227_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_227_), .Y(_228_) );
	NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_228_), .Y(reg_dataIn_13_) );
	INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_229_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(adder_result_14_), .C(_69__bF_buf0), .Y(_230_) );
	OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_71__bF_buf0), .C(_230_), .Y(_231_) );
	AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(mulOut_14_), .B(_66__bF_buf0), .C(_231_), .Y(_232_) );
	INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_14_), .Y(_233_) );
	INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_234_) );
	OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_78__bF_buf0), .C(_234_), .D(_77__bF_buf0), .Y(_235_) );
	INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_236_) );
	INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(divideOut_14_), .Y(_237_) );
	OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_83__bF_buf0), .C(_237_), .D(_82__bF_buf0), .Y(_238_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_238_), .Y(_239_) );
	NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_239_), .Y(reg_dataIn_14_) );
	INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_240_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(adder_result_15_), .C(_69__bF_buf4), .Y(_241_) );
	OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_71__bF_buf4), .C(_241_), .Y(_242_) );
	AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(mulOut_15_), .B(_66__bF_buf4), .C(_242_), .Y(_243_) );
	INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_15_), .Y(_244_) );
	INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_245_) );
	OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_78__bF_buf4), .C(_245_), .D(_77__bF_buf4), .Y(_246_) );
	INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_247_) );
	INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(divideOut_15_), .Y(_248_) );
	OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_83__bF_buf4), .C(_248_), .D(_82__bF_buf4), .Y(_249_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_249_), .Y(_250_) );
	NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_250_), .Y(reg_dataIn_15_) );
	INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_251_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_16_), .C(_69__bF_buf3), .Y(_252_) );
	OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_71__bF_buf3), .C(_252_), .Y(_253_) );
	AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(mulOut_16_), .B(_66__bF_buf3), .C(_253_), .Y(_254_) );
	INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_16_), .Y(_255_) );
	INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_256_) );
	OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_78__bF_buf3), .C(_256_), .D(_77__bF_buf3), .Y(_257_) );
	INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_258_) );
	INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(divideOut_16_), .Y(_259_) );
	OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_83__bF_buf3), .C(_259_), .D(_82__bF_buf3), .Y(_260_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_260_), .Y(_261_) );
	NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_261_), .Y(reg_dataIn_16_) );
	INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_262_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(adder_result_17_), .C(_69__bF_buf2), .Y(_263_) );
	OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_71__bF_buf2), .C(_263_), .Y(_264_) );
	AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(mulOut_17_), .B(_66__bF_buf2), .C(_264_), .Y(_265_) );
	INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_17_), .Y(_266_) );
	INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_267_) );
	OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_78__bF_buf2), .C(_267_), .D(_77__bF_buf2), .Y(_268_) );
	INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_269_) );
	INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(divideOut_17_), .Y(_270_) );
	OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_83__bF_buf2), .C(_270_), .D(_82__bF_buf2), .Y(_271_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_271_), .Y(_272_) );
	NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_272_), .Y(reg_dataIn_17_) );
	INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_273_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_18_), .C(_69__bF_buf1), .Y(_274_) );
	OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_71__bF_buf1), .C(_274_), .Y(_275_) );
	AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(mulOut_18_), .B(_66__bF_buf1), .C(_275_), .Y(_276_) );
	INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_18_), .Y(_277_) );
	INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_278_) );
	OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_78__bF_buf1), .C(_278_), .D(_77__bF_buf1), .Y(_279_) );
	INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_280_) );
	INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(divideOut_18_), .Y(_281_) );
	OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_83__bF_buf1), .C(_281_), .D(_82__bF_buf1), .Y(_282_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_282_), .Y(_283_) );
	NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_283_), .Y(reg_dataIn_18_) );
	INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_284_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(adder_result_19_), .C(_69__bF_buf0), .Y(_285_) );
	OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_71__bF_buf0), .C(_285_), .Y(_286_) );
	AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(mulOut_19_), .B(_66__bF_buf0), .C(_286_), .Y(_287_) );
	INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_19_), .Y(_288_) );
	INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_289_) );
	OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_78__bF_buf0), .C(_289_), .D(_77__bF_buf0), .Y(_290_) );
	INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_291_) );
	INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(divideOut_19_), .Y(_292_) );
	OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_83__bF_buf0), .C(_292_), .D(_82__bF_buf0), .Y(_293_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_293_), .Y(_294_) );
	NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_294_), .Y(reg_dataIn_19_) );
	INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_295_) );
	NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(adder_result_20_), .C(_69__bF_buf4), .Y(_296_) );
	OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_71__bF_buf4), .C(_296_), .Y(_297_) );
	AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(mulOut_20_), .B(_66__bF_buf4), .C(_297_), .Y(_298_) );
	INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_20_), .Y(_299_) );
	INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_300_) );
	OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_78__bF_buf4), .C(_300_), .D(_77__bF_buf4), .Y(_301_) );
	INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_302_) );
	INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(divideOut_20_), .Y(_303_) );
	OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_83__bF_buf4), .C(_303_), .D(_82__bF_buf4), .Y(_304_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_304_), .Y(_305_) );
	NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_305_), .Y(reg_dataIn_20_) );
	INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_306_) );
	NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_21_), .C(_69__bF_buf3), .Y(_307_) );
	OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_71__bF_buf3), .C(_307_), .Y(_308_) );
	AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(mulOut_21_), .B(_66__bF_buf3), .C(_308_), .Y(_309_) );
	INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_21_), .Y(_310_) );
	INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_311_) );
	OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_78__bF_buf3), .C(_311_), .D(_77__bF_buf3), .Y(_312_) );
	INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_313_) );
	INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(divideOut_21_), .Y(_314_) );
	OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_83__bF_buf3), .C(_314_), .D(_82__bF_buf3), .Y(_315_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_315_), .Y(_316_) );
	NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_316_), .Y(reg_dataIn_21_) );
	INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_317_) );
	NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(adder_result_22_), .C(_69__bF_buf2), .Y(_318_) );
	OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_71__bF_buf2), .C(_318_), .Y(_319_) );
	AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(mulOut_22_), .B(_66__bF_buf2), .C(_319_), .Y(_320_) );
	INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_22_), .Y(_321_) );
	INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_322_) );
	OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_78__bF_buf2), .C(_322_), .D(_77__bF_buf2), .Y(_323_) );
	INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_324_) );
	INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(divideOut_22_), .Y(_325_) );
	OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_83__bF_buf2), .C(_325_), .D(_82__bF_buf2), .Y(_326_) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_326_), .Y(_327_) );
	NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_327_), .Y(reg_dataIn_22_) );
	INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_328_) );
	NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_23_), .C(_69__bF_buf1), .Y(_329_) );
	OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_71__bF_buf1), .C(_329_), .Y(_330_) );
	AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(mulOut_23_), .B(_66__bF_buf1), .C(_330_), .Y(_331_) );
	INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_23_), .Y(_332_) );
	INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_333_) );
	OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_78__bF_buf1), .C(_333_), .D(_77__bF_buf1), .Y(_334_) );
	INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_335_) );
	INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(divideOut_23_), .Y(_336_) );
	OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_83__bF_buf1), .C(_336_), .D(_82__bF_buf1), .Y(_337_) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_337_), .Y(_338_) );
	NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_338_), .Y(reg_dataIn_23_) );
	INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_339_) );
	NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(adder_result_24_), .C(_69__bF_buf0), .Y(_340_) );
	OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_71__bF_buf0), .C(_340_), .Y(_341_) );
	AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(mulOut_24_), .B(_66__bF_buf0), .C(_341_), .Y(_342_) );
	INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_24_), .Y(_343_) );
	INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_344_) );
	OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_78__bF_buf0), .C(_344_), .D(_77__bF_buf0), .Y(_345_) );
	INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_346_) );
	INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(divideOut_24_), .Y(_347_) );
	OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_83__bF_buf0), .C(_347_), .D(_82__bF_buf0), .Y(_348_) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_348_), .Y(_349_) );
	NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_349_), .Y(reg_dataIn_24_) );
	INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_350_) );
	NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(adder_result_25_), .C(_69__bF_buf4), .Y(_351_) );
	OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_71__bF_buf4), .C(_351_), .Y(_352_) );
	AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(mulOut_25_), .B(_66__bF_buf4), .C(_352_), .Y(_353_) );
	INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_25_), .Y(_354_) );
	INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_355_) );
	OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_78__bF_buf4), .C(_355_), .D(_77__bF_buf4), .Y(_356_) );
	INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_357_) );
	INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(divideOut_25_), .Y(_358_) );
	OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_83__bF_buf4), .C(_358_), .D(_82__bF_buf4), .Y(_359_) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_359_), .Y(_360_) );
	NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_360_), .Y(reg_dataIn_25_) );
	INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_361_) );
	NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_26_), .C(_69__bF_buf3), .Y(_362_) );
	OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_71__bF_buf3), .C(_362_), .Y(_363_) );
	AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(mulOut_26_), .B(_66__bF_buf3), .C(_363_), .Y(_364_) );
	INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_26_), .Y(_365_) );
	INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_366_) );
	OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_78__bF_buf3), .C(_366_), .D(_77__bF_buf3), .Y(_367_) );
	INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_368_) );
	INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(divideOut_26_), .Y(_369_) );
	OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_83__bF_buf3), .C(_369_), .D(_82__bF_buf3), .Y(_370_) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_370_), .Y(_371_) );
	NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_371_), .Y(reg_dataIn_26_) );
	INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_372_) );
	NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(adder_result_27_), .C(_69__bF_buf2), .Y(_373_) );
	OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_71__bF_buf2), .C(_373_), .Y(_374_) );
	AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(mulOut_27_), .B(_66__bF_buf2), .C(_374_), .Y(_375_) );
	INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_27_), .Y(_376_) );
	INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_377_) );
	OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_78__bF_buf2), .C(_377_), .D(_77__bF_buf2), .Y(_378_) );
	INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_379_) );
	INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(divideOut_27_), .Y(_380_) );
	OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_83__bF_buf2), .C(_380_), .D(_82__bF_buf2), .Y(_381_) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_381_), .Y(_382_) );
	NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_382_), .Y(reg_dataIn_27_) );
	INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_383_) );
	NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf4), .B(adder_result_28_), .C(_69__bF_buf1), .Y(_384_) );
	OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_71__bF_buf1), .C(_384_), .Y(_385_) );
	AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(mulOut_28_), .B(_66__bF_buf1), .C(_385_), .Y(_386_) );
	INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_28_), .Y(_387_) );
	INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_388_) );
	OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_78__bF_buf1), .C(_388_), .D(_77__bF_buf1), .Y(_389_) );
	INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_390_) );
	INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(divideOut_28_), .Y(_391_) );
	OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_83__bF_buf1), .C(_391_), .D(_82__bF_buf1), .Y(_392_) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_392_), .Y(_393_) );
	NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_393_), .Y(reg_dataIn_28_) );
	INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_394_) );
	NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(adder_result_29_), .C(_69__bF_buf0), .Y(_395_) );
	OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_71__bF_buf0), .C(_395_), .Y(_396_) );
	AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(mulOut_29_), .B(_66__bF_buf0), .C(_396_), .Y(_397_) );
	INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_29_), .Y(_398_) );
	INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_399_) );
	OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_78__bF_buf0), .C(_399_), .D(_77__bF_buf0), .Y(_400_) );
	INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_401_) );
	INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(divideOut_29_), .Y(_402_) );
	OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_83__bF_buf0), .C(_402_), .D(_82__bF_buf0), .Y(_403_) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_403_), .Y(_404_) );
	NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_404_), .Y(reg_dataIn_29_) );
	INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_405_) );
	NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(adder_result_30_), .C(_69__bF_buf4), .Y(_406_) );
	OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_71__bF_buf4), .C(_406_), .Y(_407_) );
	AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(mulOut_30_), .B(_66__bF_buf4), .C(_407_), .Y(_408_) );
	INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_30_), .Y(_409_) );
	INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_410_) );
	OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_78__bF_buf4), .C(_410_), .D(_77__bF_buf4), .Y(_411_) );
	INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_412_) );
	INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(divideOut_30_), .Y(_413_) );
	OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_83__bF_buf4), .C(_413_), .D(_82__bF_buf4), .Y(_414_) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_414_), .Y(_415_) );
	NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_415_), .Y(reg_dataIn_30_) );
	INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_416_) );
	NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(adder_result_31_), .C(_69__bF_buf3), .Y(_417_) );
	OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_71__bF_buf3), .C(_417_), .Y(_418_) );
	AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(mulOut_31_), .B(_66__bF_buf3), .C(_418_), .Y(_419_) );
	INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_result_31_), .Y(_420_) );
	INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_421_) );
	OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_78__bF_buf3), .C(_421_), .D(_77__bF_buf3), .Y(_422_) );
	INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_423_) );
	INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(divideOut_31_), .Y(_424_) );
	OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_83__bF_buf3), .C(_424_), .D(_82__bF_buf3), .Y(_425_) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_425_), .Y(_426_) );
	NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_426_), .Y(reg_dataIn_31_) );
	BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(_427_), .Y(busy) );
	BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(_428__0_), .Y(tempRegOut[0]) );
	BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(_428__1_), .Y(tempRegOut[1]) );
	BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(_428__2_), .Y(tempRegOut[2]) );
	BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(_428__3_), .Y(tempRegOut[3]) );
	BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(_428__4_), .Y(tempRegOut[4]) );
	BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(_428__5_), .Y(tempRegOut[5]) );
	BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(_428__6_), .Y(tempRegOut[6]) );
	BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(_428__7_), .Y(tempRegOut[7]) );
	BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(_428__8_), .Y(tempRegOut[8]) );
	BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(_428__9_), .Y(tempRegOut[9]) );
	BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(_428__10_), .Y(tempRegOut[10]) );
	BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(_428__11_), .Y(tempRegOut[11]) );
	BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(_428__12_), .Y(tempRegOut[12]) );
	BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(_428__13_), .Y(tempRegOut[13]) );
	BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(_428__14_), .Y(tempRegOut[14]) );
	BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(_428__15_), .Y(tempRegOut[15]) );
	BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(_428__16_), .Y(tempRegOut[16]) );
	BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(_428__17_), .Y(tempRegOut[17]) );
	BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(_428__18_), .Y(tempRegOut[18]) );
	BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(_428__19_), .Y(tempRegOut[19]) );
	BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(_428__20_), .Y(tempRegOut[20]) );
	BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(_428__21_), .Y(tempRegOut[21]) );
	BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(_428__22_), .Y(tempRegOut[22]) );
	BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(_428__23_), .Y(tempRegOut[23]) );
	BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(_428__24_), .Y(tempRegOut[24]) );
	BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(_428__25_), .Y(tempRegOut[25]) );
	BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(_428__26_), .Y(tempRegOut[26]) );
	BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(_428__27_), .Y(tempRegOut[27]) );
	BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(_428__28_), .Y(tempRegOut[28]) );
	BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(_428__29_), .Y(tempRegOut[29]) );
	BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(_428__30_), .Y(tempRegOut[30]) );
	BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(_428__31_), .Y(tempRegOut[31]) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf4), .B(adder_bOperand_0_bF_buf6), .Y(adder_result_0_) );
	XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf5), .B(adder_bOperand_1_bF_buf6), .Y(_914_) );
	INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf3), .Y(_429_) );
	INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .Y(_430_) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_430_), .Y(_431_) );
	OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf2), .B(_430_), .C(adder_subtract_bF_buf3), .Y(_432_) );
	OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf2), .B(_431_), .C(_432_), .Y(_433_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_914_), .Y(adder_result_1_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf4), .B(adder_bOperand_2_bF_buf5), .Y(_434_) );
	INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf1), .Y(_435_) );
	INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf4), .Y(_436_) );
	INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .Y(_437_) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_437_), .Y(_438_) );
	AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_431_), .C(_438_), .Y(_439_) );
	OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf1), .B(_430_), .C(aOperand_frameOut_1_bF_buf3), .D(_437_), .Y(_440_) );
	OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(adder_bOperand_1_bF_buf4), .C(_440_), .Y(_441_) );
	MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_441_), .S(_435__bF_buf5), .Y(_442_) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_434_), .Y(adder_result_2_) );
	INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf4), .Y(_443_) );
	NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf5), .B(_443_), .Y(_444_) );
	INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .Y(_445_) );
	NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf3), .B(_445_), .Y(_446_) );
	NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_446_), .Y(_447_) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_439_), .Y(_448_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf3), .Y(_449_) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .B(_449_), .Y(_450_) );
	NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf2), .B(_437_), .Y(_451_) );
	XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf2), .B(adder_bOperand_2_bF_buf3), .Y(_452_) );
	AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_440_), .C(_452_), .Y(_453_) );
	OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_453_), .C(adder_subtract_bF_buf0), .Y(_454_) );
	INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf2), .Y(_455_) );
	OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_455_), .C(_435__bF_buf4), .Y(_456_) );
	OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_448_), .C(_454_), .Y(_457_) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_447_), .Y(adder_result_3_) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf4), .B(adder_bOperand_4_bF_buf5), .Y(_458_) );
	NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_455_), .Y(_459_) );
	NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_445_), .Y(_460_) );
	AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_459_), .C(_460_), .Y(_461_) );
	NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_447_), .Y(_462_) );
	OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_439_), .C(_461_), .Y(_463_) );
	NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf3), .B(_463_), .Y(_464_) );
	INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_451_), .Y(_465_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(adder_bOperand_0_bF_buf4), .C(_436_), .D(adder_bOperand_1_bF_buf3), .Y(_466_) );
	OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_465_), .C(_434_), .Y(_467_) );
	OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(adder_bOperand_2_bF_buf1), .C(_446_), .Y(_468_) );
	INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_468_), .Y(_469_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(adder_bOperand_3_bF_buf3), .C(_469_), .D(_467_), .Y(_470_) );
	OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_470_), .C(_464_), .Y(_471_) );
	XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_458_), .Y(adder_result_4_) );
	INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf4), .Y(_472_) );
	NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf4), .B(_472_), .Y(_473_) );
	INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf3), .Y(_474_) );
	NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf3), .B(_474_), .Y(_475_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_475_), .Y(_476_) );
	INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .Y(_477_) );
	NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .B(_477_), .Y(_478_) );
	INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf2), .Y(_479_) );
	NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf3), .B(_479_), .Y(_480_) );
	NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_478_), .Y(_481_) );
	OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_453_), .C(_444_), .Y(_482_) );
	OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_482_), .C(_478_), .Y(_483_) );
	INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_463_), .Y(_484_) );
	NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_484_), .Y(_485_) );
	NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_477_), .Y(_486_) );
	OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_485_), .C(_435__bF_buf1), .Y(_487_) );
	OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf0), .B(_483_), .C(_487_), .Y(_488_) );
	XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_476_), .Y(adder_result_5_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf4), .Y(_489_) );
	NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(_489_), .Y(_490_) );
	INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf4), .Y(_491_) );
	NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf3), .B(_491_), .Y(_492_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_492_), .Y(_493_) );
	NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_476_), .Y(_494_) );
	OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(adder_bOperand_5_bF_buf2), .C(_478_), .Y(_495_) );
	OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf2), .B(_474_), .C(_495_), .Y(_496_) );
	OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_482_), .C(_496_), .Y(_497_) );
	NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_475_), .Y(_498_) );
	NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_474_), .Y(_499_) );
	AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_486_), .C(_499_), .Y(_500_) );
	NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_498_), .Y(_501_) );
	OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_484_), .C(_500_), .Y(_502_) );
	NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf5), .B(_502_), .Y(_503_) );
	OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf4), .B(_497_), .C(_503_), .Y(_504_) );
	XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_493_), .Y(adder_result_6_) );
	INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf4), .Y(_505_) );
	NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(_505_), .Y(_506_) );
	INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf4), .Y(_507_) );
	NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf3), .B(_507_), .Y(_508_) );
	NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_508_), .Y(_509_) );
	NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf3), .B(_489_), .Y(_510_) );
	OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_497_), .C(_490_), .Y(_511_) );
	NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_492_), .Y(_512_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_512_), .Y(_513_) );
	OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_491_), .C(_435__bF_buf3), .Y(_514_) );
	OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_511_), .C(_514_), .D(_513_), .Y(_515_) );
	XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_509_), .Y(adder_result_7_) );
	INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf4), .Y(_516_) );
	NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf4), .B(_516_), .Y(_517_) );
	INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf3), .Y(_518_) );
	NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf3), .B(_518_), .Y(_519_) );
	NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_519_), .Y(_520_) );
	INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_520_), .Y(_521_) );
	NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_498_), .Y(_522_) );
	NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_509_), .Y(_523_) );
	NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_523_), .Y(_524_) );
	INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(_473_), .Y(_525_) );
	OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_525_), .C(_475_), .Y(_526_) );
	OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf2), .B(_507_), .C(_510_), .Y(_527_) );
	OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(adder_bOperand_7_bF_buf3), .C(_527_), .Y(_528_) );
	AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_526_), .C(_528_), .Y(_529_) );
	OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_482_), .C(_529_), .Y(_530_) );
	NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_509_), .Y(_531_) );
	NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_531_), .Y(_532_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_532_), .Y(_533_) );
	NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_491_), .Y(_534_) );
	NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_507_), .Y(_535_) );
	AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_534_), .C(_535_), .Y(_536_) );
	OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_500_), .C(_536_), .Y(_537_) );
	OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_533_), .C(_435__bF_buf1), .Y(_538_) );
	OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf0), .B(_530_), .C(_538_), .Y(_539_) );
	XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_521_), .Y(adder_result_8_) );
	INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf4), .Y(_540_) );
	NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf4), .B(_540_), .Y(_541_) );
	INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf3), .Y(_542_) );
	NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf3), .B(_542_), .Y(_543_) );
	NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_543_), .Y(_544_) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_508_), .Y(_545_) );
	NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_545_), .Y(_546_) );
	NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_546_), .Y(_547_) );
	AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_508_), .Y(_548_) );
	OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_546_), .C(_548_), .Y(_549_) );
	AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_470_), .C(_549_), .Y(_550_) );
	OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(adder_bOperand_8_bF_buf2), .C(_550_), .Y(_551_) );
	OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf2), .B(_518_), .C(_551_), .Y(_552_) );
	AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_532_), .C(_537_), .Y(_553_) );
	NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_553_), .Y(_554_) );
	OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_518_), .C(_435__bF_buf5), .Y(_555_) );
	OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_555_), .C(_435__bF_buf4), .D(_552_), .Y(_556_) );
	XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_544_), .Y(adder_result_9_) );
	INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf4), .Y(_557_) );
	NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf4), .B(_557_), .Y(_558_) );
	INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf3), .Y(_559_) );
	NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf3), .B(_559_), .Y(_560_) );
	NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_560_), .Y(_561_) );
	NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_544_), .Y(_562_) );
	INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_541_), .Y(_563_) );
	OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_563_), .C(_543_), .Y(_564_) );
	AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_562_), .C(_564_), .Y(_565_) );
	NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf3), .B(_565_), .Y(_566_) );
	NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_518_), .Y(_567_) );
	NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .Y(_568_) );
	AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_567_), .C(_568_), .Y(_569_) );
	NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_544_), .Y(_570_) );
	OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_553_), .C(_569_), .Y(_571_) );
	INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_571_), .Y(_572_) );
	OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf2), .B(_572_), .C(_566_), .Y(_573_) );
	XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_561_), .Y(adder_result_10_) );
	INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf4), .Y(_574_) );
	NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf3), .B(_574_), .Y(_575_) );
	INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf2), .Y(_576_) );
	NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf3), .B(_576_), .Y(_577_) );
	NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_577_), .Y(_578_) );
	OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(adder_bOperand_10_bF_buf2), .C(_565_), .Y(_579_) );
	OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf2), .B(_557_), .C(_579_), .Y(_580_) );
	NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_572_), .Y(_581_) );
	OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_557_), .C(_435__bF_buf3), .Y(_582_) );
	OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_580_), .C(_582_), .D(_581_), .Y(_583_) );
	XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_578_), .Y(adder_result_11_) );
	INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf4), .Y(_584_) );
	NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf3), .B(_584_), .Y(_585_) );
	INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf2), .Y(_586_) );
	NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf3), .B(_586_), .Y(_587_) );
	AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_587_), .Y(_588_) );
	OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(adder_bOperand_9_bF_buf2), .C(_519_), .Y(_589_) );
	OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf2), .B(_542_), .C(_589_), .Y(_590_) );
	XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf1), .B(adder_bOperand_10_bF_buf1), .Y(_591_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_591_), .Y(_592_) );
	OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf2), .B(_576_), .C(_560_), .Y(_593_) );
	AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_577_), .Y(_594_) );
	OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_592_), .C(_594_), .Y(_595_) );
	NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_578_), .Y(_596_) );
	AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_596_), .Y(_597_) );
	AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_597_), .C(_595_), .Y(_598_) );
	NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf1), .B(_598_), .Y(_599_) );
	OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_560_), .C(_578_), .Y(_600_) );
	NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_557_), .Y(_601_) );
	NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_576_), .Y(_602_) );
	AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_601_), .C(_602_), .Y(_603_) );
	OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_569_), .C(_603_), .Y(_604_) );
	INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_604_), .Y(_605_) );
	NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_600_), .Y(_606_) );
	OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_533_), .C(_606_), .Y(_607_) );
	AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_605_), .Y(_608_) );
	OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf0), .B(_608_), .C(_599_), .Y(_609_) );
	XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_588_), .Y(adder_result_12_) );
	INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf4), .Y(_610_) );
	NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf3), .B(_610_), .Y(_611_) );
	INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf2), .Y(_612_) );
	NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf3), .B(_612_), .Y(_613_) );
	NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_613_), .Y(_614_) );
	OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(adder_bOperand_12_bF_buf1), .C(_598_), .Y(_615_) );
	OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf2), .B(_586_), .C(_615_), .Y(_616_) );
	NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_608_), .Y(_617_) );
	OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_586_), .C(_435__bF_buf1), .Y(_618_) );
	OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf0), .B(_616_), .C(_618_), .D(_617_), .Y(_619_) );
	XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_614_), .Y(adder_result_13_) );
	INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf4), .Y(_620_) );
	NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf3), .B(_620_), .Y(_621_) );
	INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf2), .Y(_622_) );
	NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf3), .B(_622_), .Y(_623_) );
	AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_623_), .Y(_624_) );
	AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_613_), .Y(_625_) );
	NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_625_), .Y(_626_) );
	OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(adder_bOperand_13_bF_buf1), .C(_587_), .Y(_627_) );
	OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf2), .B(_612_), .C(_627_), .Y(_628_) );
	OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_598_), .C(_628_), .Y(_629_) );
	NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_586_), .Y(_630_) );
	NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_612_), .Y(_631_) );
	AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_630_), .C(_631_), .Y(_632_) );
	INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_632_), .Y(_633_) );
	NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_587_), .Y(_634_) );
	NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_614_), .Y(_635_) );
	NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_608_), .Y(_636_) );
	OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_636_), .C(_435__bF_buf5), .Y(_637_) );
	OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf4), .B(_629_), .C(_637_), .Y(_638_) );
	XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_624_), .Y(adder_result_14_) );
	INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf4), .Y(_639_) );
	NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf4), .B(_639_), .Y(_640_) );
	INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf3), .Y(_641_) );
	NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf3), .B(_641_), .Y(_642_) );
	NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_642_), .Y(_643_) );
	NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf1), .B(_620_), .Y(_644_) );
	OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_629_), .C(_621_), .Y(_645_) );
	NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_636_), .Y(_646_) );
	NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_646_), .Y(_647_) );
	OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_622_), .C(_435__bF_buf3), .Y(_648_) );
	OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_645_), .C(_648_), .D(_647_), .Y(_649_) );
	XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_643_), .Y(adder_result_15_) );
	AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf4), .B(adder_bOperand_16_bF_buf3), .Y(_650_) );
	NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf3), .B(adder_bOperand_16_bF_buf2), .Y(_651_) );
	NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_650_), .Y(_652_) );
	INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_652_), .Y(_653_) );
	NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_623_), .Y(_654_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_643_), .Y(_655_) );
	NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_655_), .Y(_656_) );
	NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_656_), .Y(_657_) );
	OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf2), .B(_641_), .C(_644_), .Y(_658_) );
	OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(adder_bOperand_15_bF_buf2), .C(_658_), .Y(_659_) );
	INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_659_), .Y(_660_) );
	OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_655_), .C(_660_), .Y(_661_) );
	AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_656_), .C(_661_), .Y(_662_) );
	OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_550_), .C(_662_), .Y(_663_) );
	NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_643_), .Y(_664_) );
	NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_664_), .Y(_665_) );
	NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_665_), .Y(_666_) );
	NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_553_), .Y(_667_) );
	NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_622_), .Y(_668_) );
	NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_641_), .Y(_669_) );
	AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_668_), .C(_669_), .Y(_670_) );
	OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_632_), .C(_670_), .Y(_671_) );
	AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_665_), .C(_671_), .Y(_672_) );
	INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_672_), .Y(_673_) );
	OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_667_), .C(_435__bF_buf1), .Y(_674_) );
	OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf0), .B(_663_), .C(_674_), .Y(_675_) );
	XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_653_), .Y(adder_result_16_) );
	INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf4), .Y(_676_) );
	NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf3), .B(_676_), .Y(_677_) );
	INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf2), .Y(_678_) );
	NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf3), .B(_678_), .Y(_679_) );
	NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_679_), .Y(_680_) );
	INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_680_), .Y(_681_) );
	OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_553_), .C(_672_), .Y(_682_) );
	NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf3), .B(_651_), .Y(_683_) );
	OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_682_), .C(_683_), .Y(_684_) );
	NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_562_), .Y(_685_) );
	NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_643_), .Y(_686_) );
	NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_625_), .C(_686_), .Y(_687_) );
	NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_687_), .Y(_688_) );
	OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(adder_bOperand_11_bF_buf1), .C(_593_), .Y(_689_) );
	AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_564_), .C(_689_), .Y(_690_) );
	OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_614_), .C(_613_), .Y(_691_) );
	AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_686_), .C(_659_), .Y(_692_) );
	OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_690_), .C(_692_), .Y(_693_) );
	AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_688_), .C(_693_), .Y(_694_) );
	INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_bF_buf1), .Y(_695_) );
	NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf2), .B(_695_), .Y(_696_) );
	OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_694_), .C(_696_), .Y(_697_) );
	OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf5), .B(_697_), .C(_684_), .Y(_698_) );
	XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_681_), .Y(adder_result_17_) );
	INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf4), .Y(_699_) );
	NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf3), .B(_699_), .Y(_700_) );
	INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf2), .Y(_701_) );
	NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf3), .B(_701_), .Y(_702_) );
	NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_702_), .Y(_703_) );
	INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(_703_), .Y(_704_) );
	OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_680_), .C(_679_), .Y(_705_) );
	INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_706_) );
	OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_651_), .C(_681_), .Y(_707_) );
	OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_694_), .C(_706_), .Y(_708_) );
	NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_678_), .Y(_709_) );
	AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_650_), .C(_709_), .Y(_710_) );
	INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_710_), .Y(_711_) );
	NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_681_), .Y(_712_) );
	AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_712_), .C(_711_), .Y(_713_) );
	MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_708_), .S(_435__bF_buf4), .Y(_714_) );
	XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_704_), .Y(adder_result_18_) );
	INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf4), .Y(_715_) );
	NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf3), .B(_715_), .Y(_716_) );
	INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf2), .Y(_717_) );
	NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf3), .B(_717_), .Y(_718_) );
	NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_718_), .Y(_719_) );
	INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_702_), .Y(_720_) );
	OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_708_), .C(_700_), .Y(_721_) );
	NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_713_), .Y(_722_) );
	OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_701_), .C(_435__bF_buf3), .Y(_723_) );
	OAI22X1 OAI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_721_), .C(_723_), .D(_722_), .Y(_724_) );
	XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_719_), .Y(adder_result_19_) );
	INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf4), .Y(_725_) );
	NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf3), .B(_725_), .Y(_726_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(adder_bOperand_20_bF_buf2), .Y(_727_) );
	NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_727_), .Y(_728_) );
	INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(_728_), .Y(_729_) );
	OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_719_), .C(_718_), .Y(_730_) );
	NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_719_), .Y(_731_) );
	AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_731_), .C(_730_), .Y(_732_) );
	INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_731_), .Y(_733_) );
	NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_733_), .Y(_734_) );
	INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_734_), .Y(_735_) );
	OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_694_), .C(_732_), .Y(_736_) );
	INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(_682_), .Y(_737_) );
	NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_719_), .Y(_738_) );
	NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_710_), .Y(_739_) );
	INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_719_), .Y(_740_) );
	NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf2), .B(adder_bOperand_18_bF_buf1), .Y(_741_) );
	NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf2), .B(adder_bOperand_19_bF_buf1), .Y(_742_) );
	OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_740_), .C(_742_), .Y(_743_) );
	NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_739_), .Y(_744_) );
	NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_719_), .C(_712_), .Y(_745_) );
	OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_737_), .C(_744_), .Y(_746_) );
	NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf1), .B(_746_), .Y(_747_) );
	OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf0), .B(_736_), .C(_747_), .Y(_748_) );
	XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_729_), .Y(adder_result_20_) );
	INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf4), .Y(_749_) );
	NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf3), .B(_749_), .Y(_750_) );
	INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf2), .Y(_751_) );
	NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf3), .B(_751_), .Y(_752_) );
	NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_752_), .Y(_753_) );
	NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf3), .B(adder_bOperand_20_bF_buf1), .Y(_754_) );
	INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(_754_), .Y(_755_) );
	INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(_746_), .Y(_756_) );
	OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_756_), .C(_435__bF_buf5), .Y(_757_) );
	INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(_736_), .Y(_758_) );
	OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(adder_bOperand_20_bF_buf0), .C(_758_), .Y(_759_) );
	NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf2), .B(_726_), .C(_759_), .Y(_760_) );
	OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_757_), .C(_760_), .Y(_761_) );
	XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_753_), .Y(adder_result_21_) );
	INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf3), .Y(_762_) );
	NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf3), .B(_762_), .Y(_763_) );
	INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf2), .Y(_764_) );
	NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf2), .B(_764_), .Y(_765_) );
	NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_765_), .Y(_766_) );
	NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_728_), .Y(_767_) );
	INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_767_), .Y(_768_) );
	OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(adder_bOperand_20_bF_buf3), .C(_752_), .Y(_769_) );
	OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf2), .B(_751_), .C(_769_), .Y(_770_) );
	OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_758_), .C(_770_), .Y(_771_) );
	NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf4), .B(_771_), .Y(_772_) );
	AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_752_), .Y(_773_) );
	NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf1), .B(adder_bOperand_21_bF_buf1), .Y(_774_) );
	OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_773_), .C(_774_), .Y(_775_) );
	NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_729_), .Y(_776_) );
	AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_776_), .C(_775_), .Y(_777_) );
	NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf1), .B(_777_), .Y(_778_) );
	NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_778_), .Y(_779_) );
	XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_766_), .Y(adder_result_22_) );
	XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .B(adder_bOperand_23_), .Y(_780_) );
	NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf1), .B(adder_bOperand_22_bF_buf1), .Y(_781_) );
	INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_781_), .Y(_782_) );
	OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_777_), .C(_435__bF_buf3), .Y(_783_) );
	NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_763_), .Y(_784_) );
	OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_771_), .C(_784_), .Y(_785_) );
	OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_783_), .C(_785_), .Y(_786_) );
	XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_780_), .Y(adder_result_23_) );
	INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .Y(_787_) );
	NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf3), .B(_787_), .Y(_788_) );
	INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf2), .Y(_789_) );
	NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .B(_789_), .Y(_790_) );
	NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_790_), .Y(_791_) );
	NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_780_), .C(_767_), .Y(_792_) );
	NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_735_), .Y(_793_) );
	NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_792_), .Y(_794_) );
	NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_766_), .Y(_795_) );
	INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .Y(_796_) );
	NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_23_), .B(_796_), .Y(_797_) );
	AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_765_), .C(_797_), .Y(_798_) );
	OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_795_), .C(_798_), .Y(_799_) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_799_), .Y(_800_) );
	AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_793_), .C(_800_), .Y(_801_) );
	NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf0), .B(_801_), .Y(_802_) );
	NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_766_), .Y(_803_) );
	NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_803_), .B(_776_), .Y(_804_) );
	NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_804_), .Y(_805_) );
	NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .B(adder_bOperand_23_), .Y(_806_) );
	OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_780_), .C(_806_), .Y(_807_) );
	AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_803_), .C(_807_), .Y(_808_) );
	OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_744_), .C(_808_), .Y(_809_) );
	AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_805_), .C(_809_), .Y(_810_) );
	OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf3), .B(_810_), .C(_802_), .Y(_811_) );
	XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_791_), .Y(adder_result_24_) );
	INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf3), .Y(_812_) );
	NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_25_), .B(_812_), .Y(_813_) );
	INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_25_), .Y(_814_) );
	NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf2), .B(_814_), .Y(_815_) );
	NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_815_), .Y(_816_) );
	INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(_792_), .Y(_817_) );
	NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_817_), .Y(_818_) );
	NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_794_), .Y(_819_) );
	OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_694_), .C(_819_), .Y(_820_) );
	AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_820_), .B(_791_), .C(_790_), .Y(_821_) );
	NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_810_), .Y(_822_) );
	OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_787_), .C(_435__bF_buf1), .Y(_823_) );
	OAI22X1 OAI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf0), .B(_821_), .C(_823_), .D(_822_), .Y(_824_) );
	XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_816_), .Y(adder_result_25_) );
	INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_26_), .Y(_825_) );
	NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_26_), .B(_825_), .Y(_826_) );
	INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_26_), .Y(_827_) );
	NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_26_), .B(_827_), .Y(_828_) );
	NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_828_), .Y(_829_) );
	INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_829_), .Y(_830_) );
	INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(_816_), .Y(_831_) );
	NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_831_), .Y(_832_) );
	OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(adder_bOperand_24_), .C(_815_), .Y(_833_) );
	OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf1), .B(_814_), .C(_833_), .Y(_834_) );
	OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_801_), .C(_834_), .Y(_835_) );
	INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(_810_), .Y(_836_) );
	NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf1), .B(adder_bOperand_24_), .C(_816_), .Y(_837_) );
	OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_814_), .C(_837_), .Y(_838_) );
	OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_790_), .C(_816_), .Y(_839_) );
	INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(_839_), .Y(_840_) );
	AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_840_), .C(_838_), .Y(_841_) );
	MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_835_), .S(_435__bF_buf5), .Y(_842_) );
	XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_842_), .B(_830_), .Y(adder_result_26_) );
	INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_27_), .Y(_843_) );
	INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_27_), .Y(_844_) );
	NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_844_), .Y(_845_) );
	NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_27_), .B(adder_bOperand_27_), .Y(_846_) );
	NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_845_), .Y(_847_) );
	INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(_828_), .Y(_848_) );
	OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_835_), .C(_826_), .Y(_849_) );
	NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_841_), .Y(_850_) );
	OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_827_), .C(_435__bF_buf4), .Y(_851_) );
	OAI22X1 OAI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf3), .B(_849_), .C(_851_), .D(_850_), .Y(_852_) );
	XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_847_), .Y(adder_result_27_) );
	AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_28_), .B(adder_bOperand_28_), .Y(_853_) );
	NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_28_), .B(adder_bOperand_28_), .Y(_854_) );
	NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_853_), .Y(_855_) );
	INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(_855_), .Y(_856_) );
	OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_846_), .C(_830_), .Y(_857_) );
	NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_857_), .Y(_858_) );
	INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(_858_), .Y(_859_) );
	NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_857_), .Y(_860_) );
	OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_846_), .C(_848_), .Y(_861_) );
	OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(adder_bOperand_27_), .C(_861_), .Y(_862_) );
	NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_860_), .Y(_863_) );
	OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_801_), .C(_863_), .Y(_864_) );
	AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_829_), .Y(_865_) );
	NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_865_), .Y(_866_) );
	NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_26_), .B(adder_bOperand_26_), .C(_847_), .Y(_867_) );
	OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_844_), .C(_867_), .Y(_868_) );
	AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_838_), .C(_868_), .Y(_869_) );
	OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_810_), .C(_869_), .Y(_870_) );
	NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf2), .B(_870_), .Y(_871_) );
	OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf1), .B(_864_), .C(_871_), .Y(_872_) );
	XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_856_), .Y(adder_result_28_) );
	INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .Y(_873_) );
	INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_29_), .Y(_874_) );
	NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_874_), .Y(_875_) );
	NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .B(adder_bOperand_29_), .Y(_876_) );
	NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_875_), .Y(_877_) );
	INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_877_), .Y(_878_) );
	AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_870_), .B(_855_), .C(_853_), .Y(_879_) );
	INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(_863_), .Y(_880_) );
	AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_820_), .B(_858_), .C(_880_), .Y(_881_) );
	NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_881_), .Y(_882_) );
	INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_28_), .Y(_883_) );
	OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_28_), .B(_883_), .C(adder_subtract_bF_buf2), .Y(_884_) );
	OAI22X1 OAI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_882_), .B(_884_), .C(adder_subtract_bF_buf1), .D(_879_), .Y(_885_) );
	XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_878_), .Y(adder_result_29_) );
	NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .B(adder_bOperand_30_), .Y(_886_) );
	NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .B(adder_bOperand_30_), .Y(_887_) );
	INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(_887_), .Y(_888_) );
	NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_888_), .Y(_889_) );
	OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_876_), .C(_856_), .Y(_890_) );
	NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_28_), .B(_883_), .Y(_891_) );
	NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_29_), .B(_873_), .Y(_892_) );
	AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_891_), .C(_892_), .Y(_893_) );
	OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_890_), .B(_881_), .C(_893_), .Y(_894_) );
	NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_878_), .Y(_895_) );
	OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .B(adder_bOperand_29_), .C(_853_), .Y(_896_) );
	OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_874_), .C(_896_), .Y(_897_) );
	AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_870_), .B(_895_), .C(_897_), .Y(_898_) );
	MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_894_), .S(_435__bF_buf0), .Y(_899_) );
	XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_889_), .Y(adder_result_30_) );
	XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .B(divider_absoluteValue_B_msb), .Y(_900_) );
	AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .B(adder_bOperand_30_), .C(adder_subtract_bF_buf0), .Y(_901_) );
	OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_898_), .C(_901_), .Y(_902_) );
	INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .Y(_903_) );
	NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_30_), .B(_903_), .Y(_904_) );
	INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(_890_), .Y(_905_) );
	NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_864_), .Y(_906_) );
	AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_888_), .C(_893_), .D(_906_), .Y(_907_) );
	OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_907_), .C(adder_subtract_bF_buf3), .Y(_908_) );
	NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_902_), .C(_908_), .Y(_909_) );
	INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(_900_), .Y(_910_) );
	AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_889_), .C(_904_), .Y(_911_) );
	OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_435__bF_buf5), .B(_911_), .C(_902_), .Y(_912_) );
	NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_912_), .Y(_913_) );
	NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_913_), .Y(adder_result_31_) );
	INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .Y(_1067_) );
	INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .Y(_1068_) );
	AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .B(divider_absoluteValue_B_msb), .C(adder_bOperand_30_), .D(_1068_), .Y(_1069_) );
	INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_msb), .Y(_1070_) );
	NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .B(_1070_), .Y(_1071_) );
	OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(adder_bOperand_30_), .Y(_1072_) );
	NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1069_), .C(_1072_), .Y(_1073_) );
	XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_29_), .B(aOperand_frameOut_29_), .Y(_1074_) );
	XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_28_), .B(aOperand_frameOut_28_), .Y(_1075_) );
	NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1075_), .Y(_1076_) );
	NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1076_), .Y(_1077_) );
	INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_25_), .Y(_1078_) );
	NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf0), .B(_1078_), .Y(_1079_) );
	INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .Y(_1080_) );
	NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf3), .B(_1078_), .Y(_1081_) );
	XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .B(aOperand_frameOut_24_bF_buf0), .Y(_1082_) );
	NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_1082_), .C(_1080_), .Y(_1083_) );
	INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_27_), .Y(_1084_) );
	INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_26_), .Y(_1085_) );
	AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(adder_bOperand_27_), .C(adder_bOperand_26_), .D(_1085_), .Y(_1086_) );
	INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_27_), .Y(_1087_) );
	NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_27_), .B(_1087_), .Y(_1088_) );
	OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(adder_bOperand_26_), .Y(_1089_) );
	NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1088_), .B(_1086_), .C(_1089_), .Y(_1090_) );
	NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1083_), .Y(_1091_) );
	NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1091_), .Y(_1092_) );
	INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_23_), .Y(_1093_) );
	INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf0), .Y(_1094_) );
	NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf0), .B(_1094_), .Y(_1095_) );
	OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(aOperand_frameOut_23_), .C(_1095_), .Y(_1096_) );
	NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .B(_1093_), .Y(_1097_) );
	OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf3), .B(_1094_), .C(_1097_), .Y(_1098_) );
	NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1098_), .Y(_915_) );
	XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf0), .B(aOperand_frameOut_21_bF_buf0), .Y(_916_) );
	XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf2), .B(aOperand_frameOut_20_bF_buf2), .Y(_917_) );
	NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_916_), .Y(_918_) );
	INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(_918_), .Y(_919_) );
	INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf1), .Y(_920_) );
	INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf1), .Y(_921_) );
	AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(adder_bOperand_19_bF_buf0), .C(adder_bOperand_18_bF_buf0), .D(_921_), .Y(_922_) );
	INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf3), .Y(_923_) );
	NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf0), .B(_923_), .Y(_924_) );
	INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf3), .Y(_925_) );
	NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf0), .B(_925_), .Y(_926_) );
	NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_926_), .C(_922_), .Y(_927_) );
	INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf1), .Y(_928_) );
	NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf2), .B(_928_), .Y(_929_) );
	INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_bF_buf0), .Y(_930_) );
	OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(aOperand_frameOut_16_bF_buf1), .Y(_931_) );
	INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf1), .Y(_932_) );
	AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(adder_bOperand_17_bF_buf0), .C(_930_), .D(aOperand_frameOut_16_bF_buf0), .Y(_933_) );
	NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_933_), .C(_931_), .Y(_934_) );
	NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_934_), .Y(_935_) );
	NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_915_), .B(_919_), .C(_935_), .Y(_936_) );
	NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_1092_), .Y(_937_) );
	INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf1), .Y(_938_) );
	INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf2), .Y(_939_) );
	AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(adder_bOperand_7_bF_buf2), .C(adder_bOperand_6_bF_buf2), .D(_939_), .Y(_940_) );
	INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf1), .Y(_941_) );
	NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf0), .B(_941_), .Y(_942_) );
	INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf1), .Y(_943_) );
	NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf1), .B(_943_), .Y(_944_) );
	NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_944_), .C(_940_), .Y(_945_) );
	XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf1), .B(aOperand_frameOut_5_bF_buf1), .Y(_946_) );
	XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf2), .B(aOperand_frameOut_4_bF_buf1), .Y(_947_) );
	NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_947_), .Y(_948_) );
	NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_948_), .Y(_949_) );
	INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .Y(_950_) );
	NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf0), .B(_950_), .Y(_951_) );
	INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .Y(_952_) );
	NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf1), .B(_952_), .Y(_953_) );
	NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_953_), .Y(_954_) );
	OAI22X1 OAI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf0), .B(_952_), .C(_950_), .D(aOperand_frameOut_0_bF_buf4), .Y(_955_) );
	NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_954_), .Y(_956_) );
	INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .Y(_957_) );
	INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf1), .Y(_958_) );
	AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(adder_bOperand_3_bF_buf2), .C(adder_bOperand_2_bF_buf0), .D(_958_), .Y(_959_) );
	INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf1), .Y(_960_) );
	NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(_960_), .Y(_961_) );
	INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf5), .Y(_962_) );
	NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf0), .B(_962_), .Y(_963_) );
	NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_963_), .C(_959_), .Y(_964_) );
	INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(_964_), .Y(_965_) );
	NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_965_), .C(_949_), .Y(_966_) );
	INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf1), .Y(_967_) );
	NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf1), .B(_967_), .Y(_968_) );
	INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf0), .Y(_969_) );
	OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(aOperand_frameOut_14_bF_buf2), .Y(_970_) );
	INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf0), .Y(_971_) );
	AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(aOperand_frameOut_15_bF_buf0), .C(_969_), .D(aOperand_frameOut_14_bF_buf1), .Y(_972_) );
	NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_972_), .C(_970_), .Y(_973_) );
	INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf0), .Y(_974_) );
	OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(aOperand_frameOut_13_bF_buf1), .Y(_975_) );
	NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf0), .B(_974_), .Y(_976_) );
	XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf0), .B(aOperand_frameOut_12_bF_buf1), .Y(_977_) );
	NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_976_), .C(_977_), .Y(_978_) );
	NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_978_), .Y(_979_) );
	INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf1), .Y(_980_) );
	OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(aOperand_frameOut_9_bF_buf1), .Y(_981_) );
	NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf0), .B(_980_), .Y(_982_) );
	XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf1), .B(aOperand_frameOut_8_bF_buf1), .Y(_983_) );
	NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(_982_), .C(_983_), .Y(_984_) );
	INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf1), .Y(_985_) );
	INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf0), .Y(_986_) );
	AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(adder_bOperand_11_bF_buf0), .C(adder_bOperand_10_bF_buf0), .D(_986_), .Y(_987_) );
	OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(adder_bOperand_11_bF_buf3), .Y(_988_) );
	OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(adder_bOperand_10_bF_buf4), .Y(_989_) );
	NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_988_), .C(_989_), .Y(_990_) );
	NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_984_), .Y(_991_) );
	NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_979_), .B(_991_), .Y(_992_) );
	NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_992_), .B(_966_), .Y(_993_) );
	AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_937_), .Y(comparator_equal_0_) );
	AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_915_), .Y(_994_) );
	NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf4), .B(_930_), .Y(_995_) );
	NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf0), .B(_928_), .Y(_996_) );
	AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_995_), .B(_929_), .C(_996_), .Y(_997_) );
	OAI22X1 OAI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf4), .B(_923_), .C(_925_), .D(aOperand_frameOut_18_bF_buf4), .Y(_998_) );
	OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf2), .B(_920_), .C(_998_), .Y(_999_) );
	OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_927_), .C(_999_), .Y(_1000_) );
	INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf3), .Y(_1001_) );
	INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf1), .Y(_1002_) );
	NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf4), .B(_1001_), .Y(_1003_) );
	NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf1), .B(_1002_), .C(_1003_), .Y(_1004_) );
	OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(aOperand_frameOut_21_bF_buf3), .C(_1004_), .Y(_1005_) );
	NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_915_), .Y(_1006_) );
	NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .B(_1096_), .Y(_1007_) );
	NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_1006_), .Y(_1008_) );
	AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_1000_), .C(_1008_), .Y(_1009_) );
	INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .Y(_1010_) );
	INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_29_), .Y(_1011_) );
	NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .B(_1011_), .Y(_1012_) );
	NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .B(_1011_), .Y(_1013_) );
	INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_28_), .Y(_1014_) );
	NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_28_), .B(_1014_), .Y(_1015_) );
	AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1013_), .C(_1012_), .Y(_1016_) );
	OAI22X1 OAI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1010_), .C(_1016_), .D(_1073_), .Y(_1017_) );
	INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .Y(_1018_) );
	NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf3), .B(_1018_), .Y(_1019_) );
	AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1081_), .C(_1079_), .Y(_1020_) );
	AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(aOperand_frameOut_27_), .C(_1086_), .Y(_1021_) );
	INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .Y(_1022_) );
	OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1090_), .C(_1022_), .Y(_1023_) );
	AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1077_), .C(_1017_), .Y(_1024_) );
	OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_1009_), .C(_1024_), .Y(_1025_) );
	NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf5), .B(_952_), .Y(_1026_) );
	AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_953_), .C(_1026_), .Y(_1027_) );
	NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf0), .B(_960_), .Y(_1028_) );
	NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf4), .B(_962_), .Y(_1029_) );
	OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1029_), .C(_961_), .Y(_1030_) );
	OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_964_), .C(_1030_), .Y(_1031_) );
	INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(_942_), .Y(_1032_) );
	INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf0), .Y(_1033_) );
	NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf0), .B(_1033_), .Y(_1034_) );
	NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf4), .B(_1033_), .Y(_1035_) );
	INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf1), .Y(_1036_) );
	NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf0), .B(_1036_), .Y(_1037_) );
	AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_1035_), .C(_1034_), .Y(_1038_) );
	OAI22X1 OAI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_1032_), .C(_1038_), .D(_945_), .Y(_1039_) );
	AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_1031_), .C(_1039_), .Y(_1040_) );
	NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf4), .B(_974_), .Y(_1041_) );
	INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf3), .Y(_1042_) );
	NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf0), .B(_1042_), .Y(_1043_) );
	AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .B(_976_), .C(_1041_), .Y(_1044_) );
	OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(aOperand_frameOut_14_bF_buf0), .C(_968_), .Y(_1045_) );
	OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf4), .B(_967_), .C(_1045_), .Y(_1046_) );
	OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_973_), .C(_1046_), .Y(_1047_) );
	INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(_988_), .Y(_1048_) );
	NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf4), .B(_980_), .Y(_1049_) );
	INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf0), .Y(_1050_) );
	NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf0), .B(_1050_), .Y(_1051_) );
	AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_982_), .C(_1049_), .Y(_1052_) );
	OAI22X1 OAI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_1048_), .C(_1052_), .D(_990_), .Y(_1053_) );
	AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_979_), .C(_1047_), .Y(_1054_) );
	OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_992_), .B(_1040_), .C(_1054_), .Y(_1055_) );
	AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_1055_), .C(_1025_), .Y(comparator_greater_0_) );
	INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .Y(_1056_) );
	NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_915_), .B(_919_), .Y(_1057_) );
	INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1058_) );
	AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1097_), .C(_1005_), .D(_915_), .Y(_1059_) );
	OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1058_), .C(_1059_), .Y(_1060_) );
	INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .Y(_1061_) );
	NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1077_), .Y(_1062_) );
	AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1021_), .C(_1017_), .Y(_1063_) );
	OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1020_), .C(_1063_), .Y(_1064_) );
	AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1056_), .B(_1060_), .C(_1064_), .Y(_1065_) );
	NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_1055_), .Y(_1066_) );
	AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_993_), .C(_1065_), .D(_1066_), .Y(comparator_less_0_) );
	NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .Y(_1418_) );
	NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .Y(_1429_) );
	NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1429_), .Y(_1440_) );
	NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .B(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .Y(_1451_) );
	NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .B(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .Y(_1462_) );
	NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_1462_), .Y(_1473_) );
	NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .B(_1473_), .Y(_1483_) );
	INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .Y(_1494_) );
	INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .Y(_1505_) );
	NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .Y(_1516_) );
	NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf4), .B(_1505__bF_buf4), .C(_1516_), .Y(_1527_) );
	INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .Y(_1538_) );
	INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_30_), .Y(_1549_) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_31_), .Y(_1560_) );
	NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1549_), .C(_1560__bF_buf3), .Y(_1571_) );
	NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(divider_absoluteValue_B_flipSign_result_28_), .Y(_1582_) );
	NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(divider_absoluteValue_B_flipSign_result_26_bF_buf3), .Y(_1593_) );
	NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1582_), .B(_1593_), .Y(_1604_) );
	NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1604_), .Y(_1615_) );
	NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf3), .B(divider_absoluteValue_B_flipSign_result_22_bF_buf3), .Y(_1626_) );
	NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf3), .B(divider_absoluteValue_B_flipSign_result_24_bF_buf3), .Y(_1637_) );
	NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1626_), .B(_1637_), .Y(_1648_) );
	NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_20_bF_buf3), .Y(_1659_) );
	NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_18_bF_buf4), .Y(_1670_) );
	NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1670_), .Y(_1681_) );
	NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1681_), .Y(_1692_) );
	NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf4), .B(_1692_), .Y(_1702_) );
	NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1702_), .Y(_1713_) );
	AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(_1483_), .Y(_1724_) );
	INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .Y(_1735_) );
	INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .Y(_1746_) );
	AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_1615__bF_buf3), .Y(_1757_) );
	INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .Y(_1768_) );
	NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .Y(_1779_) );
	NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf7), .B(_1735__bF_buf7), .C(_1779_), .Y(_1790_) );
	NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1790_), .Y(_1801_) );
	AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_1483_), .Y(_1812_) );
	NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf3), .B(_1812_), .Y(_1823_) );
	OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf5), .B(_1823_), .C(divider_aOp_abs_31_), .Y(_1834_) );
	NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_1757__bF_buf2), .C(_1812_), .Y(_1845_) );
	NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf6), .B(divider_aOp_abs_31_), .C(_1845_), .Y(_1856_) );
	NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_30_), .B(_1746__bF_buf4), .Y(_1867_) );
	AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1845_), .B(divider_aOp_abs_31_), .C(_1768__bF_buf5), .Y(_1878_) );
	OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_1878_), .C(_1856_), .Y(_1889_) );
	NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .B(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .Y(_1900_) );
	NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .B(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .Y(_1921_) );
	NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .B(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .Y(_1922_) );
	NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_1922_), .Y(_1933_) );
	INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .Y(_1943_) );
	NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_1779_), .C(_1943_), .Y(_1954_) );
	NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .Y(_1965_) );
	NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .Y(_1976_) );
	AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1965_), .B(_1976_), .Y(_1987_) );
	NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf2), .B(divider_absoluteValue_B_flipSign_result_23_bF_buf2), .Y(_1998_) );
	INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .Y(_2009_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .B(divider_absoluteValue_B_flipSign_result_30_), .C(divider_absoluteValue_B_flipSign_result_31_), .Y(_2020_) );
	NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_2020_), .Y(_2031_) );
	INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf2), .Y(_2042_) );
	INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .Y(_2053_) );
	NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf2), .B(divider_absoluteValue_B_flipSign_result_27_), .Y(_2064_) );
	NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf3), .B(_2053_), .C(_2064_), .Y(_2075_) );
	NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .B(_2031_), .Y(_2086_) );
	NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1998_), .B(_2086_), .Y(_2097_) );
	NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf2), .B(divider_absoluteValue_B_flipSign_result_21_bF_buf2), .Y(_2108_) );
	NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf3), .B(divider_absoluteValue_B_flipSign_result_19_bF_buf3), .Y(_2119_) );
	NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .Y(_2130_) );
	AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_2130_), .Y(_2141_) );
	NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .B(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .Y(_2152_) );
	NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_2108_), .B(_2152_), .C(_2141_), .Y(_2163_) );
	NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2097_), .Y(_2174_) );
	NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1987_), .B(_2174_), .Y(_2185_) );
	NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_2185_), .Y(_2196_) );
	AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1889_), .B(_2196_), .C(_1834_), .Y(_2207_) );
	NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_1856_), .Y(_2218_) );
	NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2196_), .B(_2218_), .Y(_2229_) );
	INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(_2229__bF_buf4), .Y(_2240_) );
	INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_31_), .Y(_2251_) );
	NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1801_), .Y(_2262_) );
	NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf3), .B(_1702_), .C(_2262_), .Y(_2272_) );
	NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_2251_), .C(_2272_), .Y(_2283_) );
	INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_2294_) );
	OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_2251_), .B(_2272_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .Y(_2305_) );
	AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .B(_2294_), .C(_2283_), .Y(_2316_) );
	OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .B(_1954_), .Y(_2327_) );
	OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_2327_), .B(_2316_), .C(divider_aOp_abs_30_), .Y(_2338_) );
	INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_30_), .Y(_2349_) );
	NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(_2349_), .Y(_2360_) );
	NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_2360_), .Y(_2371_) );
	INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(_2371_), .Y(_2382_) );
	NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .B(_2196_), .C(_1889_), .Y(_2393_) );
	AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_2338_), .B(_2393_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .Y(_2404_) );
	NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .B(_2393_), .C(_2338_), .Y(_2415_) );
	NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_29_), .B(_1746__bF_buf2), .Y(_2426_) );
	INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .Y(_2437_) );
	AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .B(_2437_), .C(_2404_), .Y(_2448_) );
	NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_2448_), .Y(_2459_) );
	INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .Y(_2470_) );
	NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf7), .B(_1735__bF_buf6), .C(_1429_), .Y(_2481_) );
	NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1451_), .Y(_2492_) );
	NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1713_), .Y(_2503_) );
	NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_2492_), .B(_2503_), .Y(_2514_) );
	INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .Y(_2525_) );
	NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_2481_), .B(_2525_), .Y(_2536_) );
	INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .Y(_2547_) );
	NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2371_), .B(_2196_), .C(_1889_), .Y(_2557_) );
	OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_2327_), .B(_2316_), .C(_2349_), .Y(_2568_) );
	NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_2557_), .C(_2568_), .Y(_2579_) );
	NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_2393_), .C(_2338_), .Y(_2590_) );
	AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_2579_), .B(_2590_), .C(_2426_), .Y(_2601_) );
	OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .B(_2601_), .C(_2547__bF_buf7), .Y(_2612_) );
	NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_2536_), .C(_2612_), .Y(_2623_) );
	OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2207_), .B(_2240__bF_buf4), .C(_2623_), .Y(_2634_) );
	OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf3), .B(_2207_), .C(_2547__bF_buf6), .Y(_2645_) );
	INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(_1834_), .Y(_2656_) );
	OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2327_), .B(_2316_), .C(_2656_), .Y(_2667_) );
	NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_2229__bF_buf3), .C(_2667_), .Y(_2678_) );
	NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2645_), .Y(_2689_) );
	OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2689_), .B(_2448_), .C(_2645_), .Y(_2700_) );
	NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_2557_), .C(_2568_), .Y(_2711_) );
	AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_2711_), .B(_2415_), .C(_2437_), .Y(_2722_) );
	OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_2722_), .B(_2601_), .Y(_2733_) );
	NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2700_), .C(_2733_), .Y(_2744_) );
	NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_2327_), .B(_2316_), .Y(divider_divuResult_30_) );
	OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_30_), .B(divider_divuResult_30_), .C(_2557_), .Y(_2765_) );
	INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .Y(_2776_) );
	AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_2568_), .B(_2557_), .C(_1768__bF_buf2), .Y(_2787_) );
	OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_2787_), .C(_2711_), .Y(_2798_) );
	INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(_2645_), .Y(_2809_) );
	AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_2645_), .B(_2678_), .Y(_2820_) );
	AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_2798_), .B(_2820_), .C(_2809_), .Y(_2831_) );
	OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2831_), .C(_2765_), .Y(_2842_) );
	NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_2744_), .C(_2842_), .Y(_2853_) );
	INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .Y(_2864_) );
	INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(_2765_), .Y(_2875_) );
	OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2831_), .C(_2875_), .Y(_2885_) );
	NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .B(_2722_), .Y(_2896_) );
	NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2896_), .C(_2700_), .Y(_2907_) );
	NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .B(_2907_), .C(_2885_), .Y(_2918_) );
	INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_29_), .Y(_2929_) );
	NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(_2929_), .Y(_2940_) );
	NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_2940_), .Y(_2951_) );
	NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_2951_), .C(_2700_), .Y(_2962_) );
	OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2831_), .C(_2929_), .Y(_2973_) );
	NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf1), .B(_2962_), .C(_2973_), .Y(_2984_) );
	AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_2973_), .B(_2962_), .C(_1768__bF_buf0), .Y(_2995_) );
	NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_28_), .B(_1746__bF_buf1), .Y(_3006_) );
	OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .B(_2995_), .C(_2984_), .Y(_3017_) );
	AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3017_), .B(_2918_), .C(_2864_), .Y(_3028_) );
	NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .B(_3028_), .Y(_3039_) );
	NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_2918_), .Y(_3050_) );
	INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(_2951_), .Y(_3061_) );
	NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_2536_), .B(_3061_), .C(_2700_), .Y(_3072_) );
	OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2831_), .C(divider_aOp_abs_29_), .Y(_3083_) );
	AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3083_), .B(_3072_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .Y(_3094_) );
	NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .B(_3072_), .C(_3083_), .Y(_3105_) );
	INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .Y(_3116_) );
	AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .B(_3116_), .C(_3094_), .Y(_3127_) );
	OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_3050_), .B(_3127_), .C(_2853_), .Y(_3138_) );
	NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_1965_), .Y(_3149_) );
	NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_2152_), .Y(_3160_) );
	INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .Y(_3171_) );
	NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2108_), .B(_3171__bF_buf3), .Y(_3182_) );
	INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(_3182_), .Y(_3193_) );
	NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(_3193_), .Y(_3204_) );
	NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3160_), .B(_3204__bF_buf4), .Y(_3215_) );
	INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .Y(_3226_) );
	NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_3149_), .B(_3226_), .Y(_3236_) );
	INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .Y(_3257_) );
	NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(_3257_), .Y(_3258_) );
	INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .Y(_3269_) );
	AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3138_), .B(_2470__bF_buf6), .C(_3269_), .Y(_3280_) );
	AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3280_), .B(_3039_), .C(_2634_), .Y(_3291_) );
	OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_3291_), .B(_1735__bF_buf5), .Y(_3302_) );
	NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf4), .B(_3291_), .Y(_3313_) );
	NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_2634_), .Y(_3324_) );
	INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .Y(_3335_) );
	NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .B(_2634_), .Y(_3346_) );
	NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_3335_), .Y(_3357_) );
	OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3028_), .C(_3335_), .Y(_3368_) );
	NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(_3368_), .Y(_3379_) );
	NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_3050_), .B(_3127_), .Y(_3390_) );
	AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .B(_3050_), .Y(_3401_) );
	NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_3390_), .B(_3401_), .Y(_3412_) );
	NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2831_), .Y(divider_divuResult_29_) );
	OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_2875_), .B(divider_divuResult_29_), .C(_2744_), .Y(_3433_) );
	OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .B(_3138_), .C(_3346_), .Y(_3444_) );
	OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3444_), .C(_3433_), .Y(_3455_) );
	OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_3379_), .C(_3455_), .Y(_3466_) );
	NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .B(_3466_), .Y(_3477_) );
	INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .Y(_3488_) );
	NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3444_), .Y(divider_divuResult_28_) );
	OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_3390_), .B(_3401_), .C(divider_divuResult_28_), .Y(_3509_) );
	NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .B(_3455_), .C(_3509_), .Y(_3520_) );
	NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf5), .B(_3466_), .Y(_3531_) );
	NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_3531_), .Y(_3542_) );
	OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_29_), .B(divider_divuResult_29_), .C(_2962_), .Y(_3553_) );
	INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .Y(_3564_) );
	OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3444_), .C(_3564_), .Y(_3575_) );
	NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3116_), .B(_2984_), .C(_3105_), .Y(_3586_) );
	OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .B(_2995_), .C(_3006_), .Y(_3597_) );
	NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_3586_), .B(_3597_), .Y(_3607_) );
	INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(_3607_), .Y(_3618_) );
	NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(_3618_), .C(_3368_), .Y(_3629_) );
	NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_3575_), .B(_3629_), .Y(_3640_) );
	INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .Y(_3651_) );
	NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_3651_), .Y(_3662_) );
	INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_28_), .Y(_3673_) );
	NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(_3673_), .Y(_3684_) );
	NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .B(_3684_), .Y(_3695_) );
	NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3695_), .B(_3258_), .C(_3368_), .Y(_3706_) );
	OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3444_), .C(_3673_), .Y(_3717_) );
	NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf7), .B(_3717_), .C(_3706_), .Y(_3728_) );
	INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(_3695_), .Y(_3739_) );
	NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_3258_), .C(_3368_), .Y(_3750_) );
	OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3444_), .C(divider_aOp_abs_28_), .Y(_3761_) );
	NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .B(_3761_), .C(_3750_), .Y(_3772_) );
	NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_27_), .B(_1746__bF_buf0), .Y(_3783_) );
	INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .Y(_3794_) );
	NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3794_), .B(_3728_), .C(_3772_), .Y(_3805_) );
	OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_3695_), .B(_3379_), .C(_3761_), .Y(_3816_) );
	AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .B(_2547__bF_buf4), .C(_1768__bF_buf6), .D(_3816_), .Y(_3827_) );
	NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_3827_), .Y(_3838_) );
	NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3662_), .C(_3838_), .Y(_3849_) );
	NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .B(_3488_), .C(_3849_), .Y(_3860_) );
	NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_3302_), .C(_3860_), .Y(_3871_) );
	INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .Y(divider_divuResult_27_) );
	AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_3651_), .C(_3805_), .D(_3827_), .Y(_3892_) );
	AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3892_), .B(_3542_), .C(_3477_), .Y(_3903_) );
	NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .B(_3302_), .Y(_3914_) );
	OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3903_), .C(_3313_), .Y(_3925_) );
	XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_3892_), .B(_3542_), .Y(_3936_) );
	NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_3936_), .C(_3925_), .Y(_3947_) );
	NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_3466_), .B(_3871_), .Y(_3958_) );
	NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .B(_3947_), .C(_3958_), .Y(_3969_) );
	AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_3892_), .B(_3542_), .Y(_3980_) );
	NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3892_), .Y(_3991_) );
	NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .B(_3980_), .Y(_4002_) );
	NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4002_), .C(_3925_), .Y(_4012_) );
	INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(_3466_), .Y(_4023_) );
	NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_4023_), .B(_3871_), .Y(_4034_) );
	NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_4012_), .C(_4034_), .Y(_4045_) );
	NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .B(_3903_), .Y(_4056_) );
	OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .B(_3980_), .C(_1735__bF_buf2), .Y(_4067_) );
	NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4056_), .C(_4067_), .Y(_4078_) );
	NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .B(_3291_), .C(_4078_), .Y(_4089_) );
	INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .Y(_4100_) );
	AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_3903_), .B(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .Y(_4111_) );
	OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_3903_), .C(_1724_), .Y(_4122_) );
	OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_4111_), .B(_4122_), .C(_3291_), .Y(_4133_) );
	NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf7), .B(_4133_), .Y(_4144_) );
	AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_4144_), .B(_4089_), .C(_3969_), .D(_4045_), .Y(_4155_) );
	NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_3651_), .B(_3871_), .Y(_4166_) );
	NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_3640_), .Y(_4177_) );
	NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_4177_), .B(_3662_), .Y(_4188_) );
	AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_3728_), .Y(_4199_) );
	XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4199_), .B(_4188_), .Y(_4210_) );
	NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4210_), .C(_3925_), .Y(_4221_) );
	AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_4166_), .B(_4221_), .C(_2470__bF_buf4), .Y(_4232_) );
	NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_3728_), .B(_3772_), .Y(_4243_) );
	NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_4243_), .Y(_4254_) );
	NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_4254_), .Y(_4265_) );
	NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4265_), .C(_3925_), .Y(_4276_) );
	INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(_3816_), .Y(_4287_) );
	NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_3871_), .Y(_4298_) );
	NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_4276_), .C(_4298_), .Y(_4309_) );
	NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf3), .B(_4221_), .C(_4166_), .Y(_4320_) );
	AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(_4320_), .C(_4232_), .Y(_4331_) );
	NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_3947_), .C(_3958_), .Y(_4342_) );
	OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_4133_), .B(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .Y(_4353_) );
	AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_4078_), .B(_3291_), .C(_4100__bF_buf6), .Y(_4364_) );
	OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_4342_), .B(_4364_), .C(_4353_), .Y(_4375_) );
	AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_4331_), .B(_4155_), .C(_4375_), .Y(_4386_) );
	INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_27_), .Y(_4397_) );
	NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf0), .B(_4397_), .Y(_4408_) );
	NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_4408_), .Y(_4419_) );
	NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4419_), .C(_3925_), .Y(_4429_) );
	NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_4397_), .B(_3871_), .Y(_4440_) );
	NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_4440_), .Y(_4451_) );
	INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(_4419_), .Y(_4462_) );
	NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4462_), .C(_3925_), .Y(_4473_) );
	NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_27_), .B(_3871_), .Y(_4484_) );
	NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_4473_), .C(_4484_), .Y(_4495_) );
	OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf5), .B(divider_aOp_abs_26_), .C(_4495_), .Y(_4506_) );
	OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .B(_4451_), .C(_4506_), .Y(_4517_) );
	NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_3640_), .B(_3871_), .Y(_4528_) );
	OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_4210_), .C(_4528_), .Y(_4539_) );
	NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .B(_4539_), .Y(_4550_) );
	XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_4199_), .B(_4188_), .Y(_4561_) );
	OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_4561_), .C(_4166_), .Y(_4572_) );
	NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_4572_), .Y(_4583_) );
	NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3816_), .B(_3871_), .Y(_4594_) );
	INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(_4265_), .Y(_4605_) );
	NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4605_), .C(_3925_), .Y(_4616_) );
	NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .B(_4616_), .C(_4594_), .Y(_4627_) );
	NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(_4627_), .Y(_4638_) );
	AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_4550_), .B(_4583_), .C(_4638_), .Y(_4649_) );
	NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_4517_), .C(_4649_), .Y(_4660_) );
	NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_1976_), .Y(_4671_) );
	NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_3149_), .B(_4671_), .Y(_4682_) );
	NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_4682_), .B(_2174_), .Y(_4693_) );
	AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_4660_), .B(_4386_), .C(_4693_), .Y(divider_divuResult_26_) );
	INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .Y(_4714_) );
	INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(_4133_), .Y(_4725_) );
	AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_4034_), .B(_4012_), .C(_1735__bF_buf0), .Y(_4736_) );
	AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(_3947_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .Y(_4747_) );
	NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf5), .B(_4133_), .Y(_4758_) );
	AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_4078_), .B(_3291_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .Y(_4769_) );
	OAI22X1 OAI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_4758_), .B(_4769_), .C(_4736_), .D(_4747_), .Y(_4780_) );
	NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_4561_), .C(_3925_), .Y(_4791_) );
	NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_4791_), .C(_4528_), .Y(_4802_) );
	AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .B(_4616_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .Y(_4813_) );
	AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_4528_), .B(_4791_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .Y(_4824_) );
	OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .B(_4824_), .C(_4802_), .Y(_4835_) );
	AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_4034_), .B(_4012_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .Y(_4846_) );
	NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .B(_4133_), .Y(_4857_) );
	NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .B(_4133_), .Y(_4868_) );
	AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_4846_), .B(_4868_), .C(_4857_), .Y(_4879_) );
	OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_4835_), .B(_4780_), .C(_4879_), .Y(_4889_) );
	AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_4484_), .B(_4473_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .Y(_4900_) );
	NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_26_), .B(_1746__bF_buf4), .Y(_4911_) );
	INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .Y(_4922_) );
	AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_4495_), .B(_4922_), .C(_4900_), .Y(_4933_) );
	NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_4638_), .B(_4933_), .Y(_4944_) );
	AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_4802_), .B(_4320_), .Y(_4955_) );
	AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_4955_), .Y(_4966_) );
	AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(_4966_), .C(_4889_), .Y(_4977_) );
	OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_4725_), .Y(_4988_) );
	INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .Y(_4999_) );
	OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_4133_), .B(divider_divuResult_26_), .C(_2229__bF_buf2), .Y(_5010_) );
	AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(_4627_), .Y(_5021_) );
	INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_26_), .Y(_5032_) );
	AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .B(_5032_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .D(_4451_), .Y(_5043_) );
	OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_4900_), .B(_5043_), .C(_5021_), .Y(_5054_) );
	NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4155_), .Y(_5065_) );
	OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_5054_), .B(_5065_), .C(_4386_), .Y(_5076_) );
	INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .Y(_5087_) );
	AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .B(_5087_), .C(_4133_), .Y(_5098_) );
	OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf2), .B(_5098_), .C(_4999__bF_buf6), .Y(_5109_) );
	OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_4002_), .C(_3958_), .Y(_5120_) );
	INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .Y(_5131_) );
	NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_4517_), .B(_4649_), .Y(_5142_) );
	AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_3969_), .B(_4045_), .C(_4835_), .D(_5142_), .Y(_5153_) );
	NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3969_), .B(_4045_), .Y(_5164_) );
	NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .B(_4824_), .Y(_5175_) );
	OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_4638_), .B(_4933_), .C(_5175_), .Y(_5186_) );
	AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_4802_), .C(_5164_), .Y(_5197_) );
	OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_5197_), .B(_5153_), .C(divider_divuResult_26_), .Y(_5208_) );
	OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_5131_), .B(divider_divuResult_26_), .C(_5208_), .Y(_5219_) );
	OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(_5219_), .C(_5109_), .Y(_5230_) );
	OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_5010_), .C(_5230_), .Y(_5241_) );
	NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_2229__bF_buf1), .C(_4988_), .Y(_5252_) );
	AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_5252_), .B(_5109_), .Y(_5263_) );
	OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_5120_), .Y(_5274_) );
	NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .B(_5274_), .C(_5208_), .Y(_5285_) );
	NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_5164_), .B(_4802_), .C(_5186_), .Y(_5296_) );
	INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(_5164_), .Y(_5307_) );
	NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_5307_), .B(_4835_), .C(_5142_), .Y(_5318_) );
	NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_5296_), .B(_5318_), .C(divider_divuResult_26_), .Y(_5329_) );
	OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_5131_), .Y(_5339_) );
	NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf4), .B(_5339_), .C(_5329_), .Y(_5350_) );
	NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_5285_), .B(_5350_), .Y(_5361_) );
	NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_5361_), .B(_5263_), .Y(_5372_) );
	NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_5076_), .Y(_5383_) );
	OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .B(_4944_), .C(_4955_), .Y(_5394_) );
	INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .Y(_5405_) );
	NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(_5405_), .C(_5054_), .Y(_5416_) );
	AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_5394_), .B(_5416_), .C(_5383_), .Y(_5437_) );
	AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .B(_5087_), .C(_4539_), .Y(_5438_) );
	OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_5438_), .B(_5437_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .Y(_5449_) );
	NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_5416_), .B(_5394_), .Y(_5460_) );
	NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_26_), .B(_5460_), .Y(_5471_) );
	OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(divider_divuResult_26_), .C(_5471_), .Y(_5482_) );
	NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_4638_), .B(_4933_), .Y(_5493_) );
	NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_5493_), .B(_5054_), .Y(_5504_) );
	NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_5504_), .C(_5076_), .Y(_5515_) );
	OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_4265_), .C(_4594_), .Y(_5526_) );
	INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(_5526_), .Y(_5537_) );
	OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_5537_), .Y(_5548_) );
	NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_5515_), .C(_5548_), .Y(_5559_) );
	OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .B(_5482_), .C(_5559_), .Y(_5570_) );
	INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(_5438_), .Y(_5581_) );
	AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_5581_), .B(_5471_), .C(_1735__bF_buf7), .Y(_5592_) );
	NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .B(_5438_), .C(_5437_), .Y(_5603_) );
	OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_5526_), .Y(_5614_) );
	INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(_5504_), .Y(_5625_) );
	NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .B(_5087_), .C(_5625_), .Y(_5636_) );
	NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .B(_5636_), .C(_5614_), .Y(_5647_) );
	NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_5647_), .Y(_5658_) );
	NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_5592_), .B(_5603_), .C(_5658_), .Y(_5669_) );
	INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(_4451_), .Y(_5680_) );
	OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_5680_), .Y(_5691_) );
	INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(_4900_), .Y(_5702_) );
	NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_4495_), .B(_4922_), .C(_5702_), .Y(_5713_) );
	NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_5680_), .Y(_5724_) );
	NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_4451_), .Y(_5735_) );
	NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .B(_5735_), .C(_5724_), .Y(_5746_) );
	AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_5746_), .B(_5713_), .Y(_5757_) );
	NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_5076_), .C(_5757_), .Y(_5768_) );
	AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_5691_), .B(_5768_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .Y(_5779_) );
	NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_5032_), .Y(_5790_) );
	NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .B(_5790_), .Y(_5801_) );
	INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(_5801_), .Y(_5812_) );
	NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_5812_), .B(_5087_), .C(_5076_), .Y(_5822_) );
	OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(divider_aOp_abs_26_), .Y(_5833_) );
	AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_5833_), .B(_5822_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .Y(_5844_) );
	NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_5768_), .C(_5691_), .Y(_5855_) );
	AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_5844_), .B(_5855_), .C(_5779_), .Y(_5866_) );
	NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_5801_), .B(_5087_), .C(_5076_), .Y(_5877_) );
	OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_5032_), .Y(_5888_) );
	NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_5877_), .C(_5888_), .Y(_5899_) );
	OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_26_), .B(divider_divuResult_26_), .C(_5877_), .Y(_5910_) );
	NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .B(_5910_), .Y(_5921_) );
	NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_5899_), .B(_5921_), .Y(_5932_) );
	OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4977_), .C(_4451_), .Y(_5943_) );
	NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_5713_), .B(_5746_), .Y(_5954_) );
	NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_5954_), .C(_5076_), .Y(_5975_) );
	NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_5975_), .C(_5943_), .Y(_5976_) );
	NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_25_), .B(_1746__bF_buf3), .Y(_5987_) );
	INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(_5987_), .Y(_5998_) );
	NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_5998_), .B(_5976_), .C(_5855_), .Y(_6009_) );
	OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_6009_), .B(_5932_), .C(_5866_), .Y(_6030_) );
	AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_5449_), .B(_5570_), .C(_5669_), .D(_6030_), .Y(_6031_) );
	OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .B(_6031_), .C(_5241_), .Y(_6042_) );
	AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_2229__bF_buf0), .B(_4988_), .C(_2514_), .D(_6042_), .Y(_6053_) );
	OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf1), .B(_6053_), .C(_4714__bF_buf6), .Y(_6064_) );
	NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .B(_6042_), .Y(_6075_) );
	NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(_6075_), .Y(_6086_) );
	NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_2229__bF_buf4), .C(_6086_), .Y(_6097_) );
	AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_6097_), .B(_6064_), .Y(_6108_) );
	INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_24_), .Y(_6119_) );
	NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(_6119_), .Y(_6130_) );
	NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_24_), .B(_1746__bF_buf2), .Y(_6141_) );
	INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_6141_), .Y(_6152_) );
	AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(divider_aOp_abs_25_), .C(_6130_), .Y(_6163_) );
	NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .B(_5877_), .C(_5888_), .Y(_6174_) );
	NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_5822_), .C(_5833_), .Y(_6185_) );
	NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_6174_), .B(_6185_), .Y(_6196_) );
	NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_5976_), .B(_5855_), .C(_6196_), .Y(_6207_) );
	OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_6163_), .B(_6207_), .C(_5866_), .Y(_6218_) );
	NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf6), .B(_5471_), .C(_5581_), .Y(_6229_) );
	NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_5515_), .C(_5548_), .Y(_6240_) );
	NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_5636_), .C(_5614_), .Y(_6251_) );
	NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_6240_), .B(_6251_), .Y(_6262_) );
	NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_5449_), .B(_6229_), .C(_6262_), .Y(_6273_) );
	NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_6273_), .B(_5372_), .Y(_6284_) );
	AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_5252_), .B(_5230_), .C(_6284_), .D(_6218_), .Y(_6295_) );
	INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(_5372_), .Y(_6306_) );
	NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_6229_), .B(_5449_), .Y(_6316_) );
	OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_6316_), .C(_6229_), .Y(_6327_) );
	NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_25_), .B(_1746__bF_buf1), .Y(_6338_) );
	NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_6338_), .B(_5998_), .Y(_6349_) );
	OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_6349_), .B(divider_aOp_abs_24_), .Y(_6360_) );
	NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_6360_), .B(_6207_), .Y(_6371_) );
	AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_6306_), .B(_6327_), .C(_6371_), .D(_6284_), .Y(_6382_) );
	AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_6295_), .B(_6382_), .C(_2525_), .Y(divider_divuResult_25_) );
	XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_6031_), .B(_5361_), .Y(_6403_) );
	NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_6403_), .B(divider_divuResult_25_), .Y(_6414_) );
	NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_5219_), .B(_6075_), .Y(_6425_) );
	NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_6414_), .C(_6425_), .Y(_6436_) );
	XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_6031_), .B(_5361_), .Y(_6447_) );
	NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_6447_), .B(divider_divuResult_25_), .Y(_6458_) );
	INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(_5219_), .Y(_6469_) );
	NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_6469_), .B(_6075_), .Y(_6480_) );
	NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_6458_), .C(_6480_), .Y(_6491_) );
	NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .B(_6436_), .Y(_6502_) );
	NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_5482_), .B(_6075_), .Y(_6513_) );
	INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .Y(_6524_) );
	INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(_6316_), .Y(_6535_) );
	AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_5976_), .B(_5855_), .Y(_6546_) );
	NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_6196_), .B(_5998_), .C(_6546_), .Y(_6557_) );
	AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_6240_), .B(_6251_), .C(_5866_), .D(_6557_), .Y(_6568_) );
	OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .B(_6568_), .C(_6535_), .Y(_6579_) );
	NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_6262_), .B(_6030_), .Y(_6590_) );
	NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_6316_), .C(_6590_), .Y(_6601_) );
	NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_6601_), .B(_6579_), .Y(_6612_) );
	NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_6612_), .B(divider_divuResult_25_), .Y(_6623_) );
	AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_6513_), .B(_6623_), .C(_4100__bF_buf3), .Y(_6634_) );
	NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_6623_), .C(_6513_), .Y(_6645_) );
	OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_5526_), .B(divider_divuResult_26_), .C(_5515_), .Y(_6656_) );
	NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_6262_), .B(_6030_), .Y(_6667_) );
	NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_6568_), .B(_6667_), .Y(_6678_) );
	NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_2514_), .B(_6678_), .C(_6042_), .Y(_6689_) );
	OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_6656_), .B(divider_divuResult_25_), .C(_6689_), .Y(_6700_) );
	NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf5), .B(_6700_), .Y(_6711_) );
	AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_6711_), .B(_6645_), .C(_6634_), .Y(_6722_) );
	NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_6502_), .B(_6108_), .C(_6722_), .Y(_6733_) );
	INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(_6064_), .Y(_6744_) );
	OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_6469_), .B(divider_divuResult_25_), .C(_6414_), .Y(_6755_) );
	NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .B(_6755_), .Y(_6766_) );
	AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_6766_), .B(_6097_), .C(_6744_), .Y(_6777_) );
	AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_6733_), .B(_6777_), .Y(_6788_) );
	AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_6108_), .B(_6502_), .Y(_6799_) );
	INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(_5482_), .Y(_6810_) );
	NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_6810_), .B(_6075_), .Y(_6821_) );
	NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_6535_), .C(_6590_), .Y(_6832_) );
	OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .B(_6568_), .C(_6316_), .Y(_6843_) );
	NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_6843_), .Y(_6854_) );
	NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_6854_), .B(divider_divuResult_25_), .Y(_6865_) );
	NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .B(_6865_), .C(_6821_), .Y(_6876_) );
	NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_6645_), .Y(_6886_) );
	XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_6700_), .B(_1735__bF_buf4), .Y(_6897_) );
	NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_6886_), .B(_6897_), .Y(_6908_) );
	OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_5680_), .B(divider_divuResult_26_), .C(_5975_), .Y(_6919_) );
	OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_5987_), .B(_5932_), .C(_5899_), .Y(_6930_) );
	XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .B(_6546_), .Y(_6941_) );
	INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(_6941_), .Y(_6952_) );
	NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_6952_), .B(divider_divuResult_25_), .Y(_6963_) );
	OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_6919_), .B(divider_divuResult_25_), .C(_6963_), .Y(_6974_) );
	NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf7), .B(_6974_), .Y(_6985_) );
	NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_5943_), .B(_5975_), .C(_6075_), .Y(_6996_) );
	AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_6996_), .B(_6963_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .Y(_7007_) );
	XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_6196_), .B(_5987_), .Y(_7018_) );
	NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_7018_), .B(divider_divuResult_25_), .Y(_7029_) );
	INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(_5910_), .Y(_7040_) );
	NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_7040_), .B(_6075_), .Y(_7051_) );
	AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_7051_), .B(_7029_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .Y(_7062_) );
	NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .B(_6963_), .C(_6996_), .Y(_7073_) );
	AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_7062_), .B(_7073_), .C(_7007_), .Y(_7084_) );
	NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_25_), .B(_6075_), .Y(_7095_) );
	NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_6349_), .B(divider_divuResult_25_), .Y(_7106_) );
	AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_7095_), .B(_7106_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .Y(_7117_) );
	NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .B(_7106_), .C(_7095_), .Y(_7128_) );
	AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(_7128_), .C(_7117_), .Y(_7139_) );
	OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_5910_), .B(divider_divuResult_25_), .C(_7029_), .Y(_7150_) );
	OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_7150_), .C(_7073_), .Y(_7161_) );
	AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_6985_), .B(_7161_), .C(_7139_), .D(_7084_), .Y(_7172_) );
	NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_6799_), .B(_6908_), .C(_7172_), .Y(_7183_) );
	AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_7183_), .B(_6788_), .C(_3257_), .Y(divider_divuResult_24_) );
	INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .Y(_7204_) );
	OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_6086_), .B(divider_divuResult_24_bF_buf3), .C(_2229__bF_buf3), .Y(_7215_) );
	XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_7215_), .B(_7204__bF_buf5), .Y(_7226_) );
	INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(_6502_), .Y(_7237_) );
	INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_6722_), .Y(_7248_) );
	NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_7172_), .Y(_7259_) );
	AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_7259_), .B(_7248_), .C(_7237_), .Y(_7270_) );
	NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_7237_), .B(_7248_), .C(_7259_), .Y(_7281_) );
	INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(_7281_), .Y(_7292_) );
	OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_7270_), .B(_7292_), .C(divider_divuResult_24_bF_buf2), .Y(_7303_) );
	NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_6064_), .B(_6097_), .C(_6502_), .Y(_7314_) );
	OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_7248_), .C(_6777_), .Y(_7325_) );
	AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_6645_), .Y(_7336_) );
	XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_6700_), .B(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .Y(_7347_) );
	NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_7347_), .B(_7336_), .Y(_7358_) );
	NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_7358_), .Y(_7369_) );
	AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_7172_), .C(_7325_), .Y(_7380_) );
	OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_6755_), .Y(_7391_) );
	NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .B(_7391_), .C(_7303_), .Y(_7401_) );
	NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_7150_), .Y(_7412_) );
	NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_6919_), .B(_6075_), .Y(_7423_) );
	NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_6941_), .B(divider_divuResult_25_), .Y(_7434_) );
	AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_7423_), .B(_7434_), .C(_2470__bF_buf6), .Y(_7445_) );
	OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_7412_), .C(_6985_), .Y(_7456_) );
	NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_7106_), .B(_7095_), .Y(_7467_) );
	INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(_7467_), .Y(_7478_) );
	OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf0), .B(divider_aOp_abs_24_), .C(_7128_), .Y(_7489_) );
	OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .B(_7478_), .C(_7489_), .Y(_7500_) );
	INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(_6974_), .Y(_7511_) );
	OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .B(_7511_), .C(_7161_), .Y(_7522_) );
	OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_7500_), .B(_7456_), .C(_7522_), .Y(_7533_) );
	OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_7358_), .B(_7533_), .C(_7248_), .Y(_7544_) );
	NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_6502_), .B(_7544_), .Y(_7555_) );
	NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf1), .B(_7281_), .C(_7555_), .Y(_7566_) );
	OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf0), .B(_6755_), .Y(_7577_) );
	NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf5), .B(_7566_), .C(_7577_), .Y(_7588_) );
	AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_7401_), .B(_7588_), .C(_7226_), .Y(_7599_) );
	OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_5482_), .B(divider_divuResult_25_), .C(_6865_), .Y(_7610_) );
	OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_7610_), .Y(_7621_) );
	NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_7347_), .B(_7172_), .Y(_7632_) );
	NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_6711_), .B(_6886_), .C(_7632_), .Y(_7643_) );
	OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_6897_), .B(_7533_), .C(_6711_), .Y(_7654_) );
	NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_7654_), .Y(_7665_) );
	NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf3), .B(_7643_), .C(_7665_), .Y(_7676_) );
	AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_7676_), .B(_7621_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .Y(_7687_) );
	NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .B(_7621_), .C(_7676_), .Y(_7698_) );
	OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_6700_), .Y(_7709_) );
	NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_6897_), .B(_7533_), .Y(_7720_) );
	NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_7632_), .B(_7720_), .C(divider_divuResult_24_bF_buf2), .Y(_7731_) );
	AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_7731_), .B(_7709_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .Y(_7742_) );
	AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_7742_), .B(_7698_), .C(_7687_), .Y(_7753_) );
	INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(_7753_), .Y(_7764_) );
	INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(_7215_), .Y(_7775_) );
	AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7566_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .Y(_7786_) );
	OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf4), .B(_7215_), .C(_7786_), .Y(_7807_) );
	OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .B(_7775_), .C(_7807_), .Y(_7808_) );
	AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .B(_7599_), .C(_7808_), .Y(_7819_) );
	XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_7215_), .B(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .Y(_7830_) );
	AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7566_), .C(_4714__bF_buf4), .Y(_7841_) );
	AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(_7391_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .Y(_7852_) );
	OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_7841_), .B(_7852_), .C(_7830_), .Y(_7863_) );
	OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf1), .B(_7610_), .Y(_7874_) );
	NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .B(_7654_), .Y(_7885_) );
	AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_7632_), .B(_6711_), .C(_6886_), .Y(_7896_) );
	OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_7896_), .B(_7885_), .C(divider_divuResult_24_bF_buf0), .Y(_7907_) );
	NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf3), .B(_7874_), .C(_7907_), .Y(_7918_) );
	NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_7632_), .B(_7720_), .Y(_7929_) );
	NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_7929_), .B(divider_divuResult_24_bF_buf3), .Y(_7940_) );
	INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_6700_), .Y(_7951_) );
	OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_7951_), .Y(_7962_) );
	NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_7962_), .C(_7940_), .Y(_7973_) );
	NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf1), .B(_7709_), .C(_7731_), .Y(_7984_) );
	NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_7973_), .B(_7984_), .Y(_7995_) );
	NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_7918_), .B(_7698_), .C(_7995_), .Y(_8005_) );
	NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_8005_), .B(_7863_), .Y(_8016_) );
	OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_7511_), .Y(_8027_) );
	NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_7445_), .B(_7007_), .Y(_8038_) );
	NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .B(_7150_), .Y(_8049_) );
	NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_7150_), .Y(_8060_) );
	INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(_8060_), .Y(_8071_) );
	AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_8071_), .B(_8049_), .C(_7139_), .Y(_8082_) );
	OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_7062_), .B(_8082_), .C(_8038_), .Y(_8093_) );
	INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(_8038_), .Y(_8104_) );
	INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(_8049_), .Y(_8115_) );
	OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_8060_), .C(_7500_), .Y(_8126_) );
	NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8104_), .C(_8126_), .Y(_8137_) );
	NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_8137_), .B(_8093_), .Y(_8148_) );
	NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_8148_), .B(divider_divuResult_24_bF_buf2), .Y(_8159_) );
	NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_8027_), .C(_8159_), .Y(_8170_) );
	INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .Y(_8181_) );
	OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_6974_), .Y(_8192_) );
	NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_7412_), .B(_8038_), .C(_8126_), .Y(_8203_) );
	OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_7062_), .B(_8082_), .C(_8104_), .Y(_8214_) );
	NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_8203_), .B(_8214_), .Y(_8225_) );
	NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .B(divider_divuResult_24_bF_buf1), .Y(_8236_) );
	NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_8192_), .C(_8236_), .Y(_8247_) );
	NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_6799_), .Y(_8258_) );
	OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_7533_), .B(_8258_), .C(_6788_), .Y(_8269_) );
	NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_8269_), .Y(_8280_) );
	NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_8049_), .B(_8071_), .C(_7139_), .Y(_8291_) );
	NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_8291_), .B(_8126_), .Y(_8302_) );
	INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(_8302_), .Y(_8313_) );
	INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_7150_), .Y(_8324_) );
	OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_8324_), .Y(_8345_) );
	OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_8313_), .B(_8280_), .C(_8345_), .Y(_8346_) );
	NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .B(_8346_), .Y(_8357_) );
	AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_8357_), .B(_8247_), .C(_8181_), .Y(_8368_) );
	AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .B(_8247_), .Y(_8379_) );
	NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_8302_), .B(divider_divuResult_24_bF_buf0), .Y(_8390_) );
	NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_8345_), .C(_8390_), .Y(_8401_) );
	NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_8313_), .B(divider_divuResult_24_bF_buf3), .Y(_8412_) );
	OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_7150_), .Y(_8423_) );
	NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf5), .B(_8423_), .C(_8412_), .Y(_8434_) );
	NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_8401_), .B(_8434_), .Y(_8445_) );
	NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_8445_), .B(_8379_), .Y(_8456_) );
	NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf2), .B(_7467_), .Y(_8467_) );
	NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_7117_), .B(_8467_), .Y(_8478_) );
	XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_8478_), .B(_6152_), .Y(_8489_) );
	NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_8489_), .C(_8269_), .Y(_8500_) );
	OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_7467_), .B(divider_divuResult_24_bF_buf2), .C(_8500_), .Y(_8511_) );
	NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_8511_), .Y(_8522_) );
	INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_23_), .Y(_8533_) );
	NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_6130_), .B(_6141_), .Y(_8544_) );
	NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_8544_), .C(_8269_), .Y(_8555_) );
	OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_6119_), .Y(_8566_) );
	NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .B(_8555_), .C(_8566_), .Y(_8577_) );
	OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(divider_aOp_abs_24_), .Y(_8588_) );
	INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_8544_), .Y(_8599_) );
	NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_8599_), .C(_8269_), .Y(_8610_) );
	NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf1), .B(_8610_), .C(_8588_), .Y(_8621_) );
	AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(_8533_), .C(_8577_), .D(_8621_), .Y(_8632_) );
	NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf0), .B(_8555_), .C(_8566_), .Y(_8643_) );
	OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .B(_8511_), .C(_8643_), .Y(_8654_) );
	OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_8632_), .C(_8522_), .Y(_8665_) );
	OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_8456_), .B(_8665_), .C(_8368_), .Y(_8676_) );
	NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_8016_), .B(_8676_), .Y(_8687_) );
	INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .Y(_8697_) );
	NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(_8697__bF_buf3), .Y(_8708_) );
	INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .Y(_8719_) );
	AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(_7819_), .C(_8719_), .Y(divider_divuResult_23_) );
	INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(_7698_), .Y(_8740_) );
	NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .B(_8740_), .Y(_8751_) );
	NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_7995_), .B(_8751_), .C(_7599_), .Y(_8762_) );
	OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_8302_), .B(_8280_), .C(_8423_), .Y(_8773_) );
	NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf4), .B(_8773_), .Y(_8784_) );
	NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .B(_8247_), .Y(_8795_) );
	OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_8795_), .C(_8170_), .Y(_8806_) );
	AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_8401_), .B(_8434_), .C(_8795_), .Y(_8817_) );
	NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_8610_), .C(_8588_), .Y(_8828_) );
	NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(_8533_), .Y(_8839_) );
	NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_8839_), .B(_8643_), .C(_8828_), .Y(_8850_) );
	XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_8478_), .B(_6141_), .Y(_8861_) );
	NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_8861_), .C(_8269_), .Y(_8872_) );
	OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_7478_), .B(divider_divuResult_24_bF_buf1), .C(_8872_), .Y(_8883_) );
	OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_6119_), .B(divider_divuResult_24_bF_buf0), .C(_8610_), .Y(_8894_) );
	AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_8883_), .B(_2547__bF_buf6), .C(_1768__bF_buf7), .D(_8894_), .Y(_8905_) );
	AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_8511_), .C(_8850_), .D(_8905_), .Y(_8916_) );
	AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_8916_), .B(_8817_), .C(_8806_), .Y(_8927_) );
	OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_8762_), .B(_8927_), .C(_7819_), .Y(_8938_) );
	AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_8938_), .B(_8708_), .C(_7775_), .Y(_8949_) );
	OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf0), .B(_8949_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .Y(_8960_) );
	INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .Y(_8971_) );
	NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_7775_), .Y(_8982_) );
	AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_7830_), .B(_7786_), .C(_8982_), .Y(_8993_) );
	OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_7753_), .B(_7863_), .C(_8993_), .Y(_9004_) );
	AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_8676_), .B(_8016_), .C(_9004_), .Y(_9015_) );
	OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_7215_), .Y(_9026_) );
	NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf6), .B(_2229__bF_buf2), .C(_9026_), .Y(_9037_) );
	NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_7588_), .B(_7401_), .Y(_9048_) );
	INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(_9048_), .Y(_9059_) );
	INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(_8005_), .Y(_9070_) );
	NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_9070_), .B(_8676_), .Y(_9081_) );
	AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_9081_), .B(_7753_), .C(_9059_), .Y(_9092_) );
	NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_8817_), .B(_8916_), .Y(_9103_) );
	AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_9103_), .B(_8368_), .C(_8005_), .Y(_9114_) );
	NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_9048_), .B(_7764_), .C(_9114_), .Y(_9125_) );
	OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_9092_), .B(_9125_), .C(divider_divuResult_23_), .Y(_9136_) );
	NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_8938_), .Y(_9147_) );
	NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_7566_), .B(_7577_), .C(_9147_), .Y(_9158_) );
	NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_9158_), .C(_9136_), .Y(_9169_) );
	NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(_7391_), .C(_9147_), .Y(_9180_) );
	OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_7764_), .B(_9114_), .C(_9048_), .Y(_9191_) );
	NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_7753_), .C(_9081_), .Y(_9202_) );
	NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_9202_), .B(_9191_), .C(divider_divuResult_23_), .Y(_9213_) );
	NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_9180_), .C(_9213_), .Y(_9224_) );
	AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_8960_), .B(_9037_), .C(_9224_), .D(_9169_), .Y(_9234_) );
	NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .B(_7676_), .C(_9147_), .Y(_9245_) );
	INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(_7742_), .Y(_9256_) );
	NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_7995_), .B(_8676_), .Y(_9267_) );
	NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_9256_), .B(_8751_), .C(_9267_), .Y(_9278_) );
	INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(_7995_), .Y(_9289_) );
	OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_8927_), .C(_9256_), .Y(_9300_) );
	OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .B(_8740_), .C(_9300_), .Y(_9311_) );
	NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_9278_), .B(_9311_), .C(divider_divuResult_23_), .Y(_9322_) );
	NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(_9245_), .C(_9322_), .Y(_9333_) );
	NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_7874_), .B(_7907_), .C(_9147_), .Y(_9344_) );
	NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_8751_), .B(_9300_), .Y(_9355_) );
	AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_8676_), .B(_7995_), .C(_7742_), .Y(_9366_) );
	OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_7687_), .B(_8740_), .C(_9366_), .Y(_9377_) );
	NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_9355_), .B(divider_divuResult_23_), .C(_9377_), .Y(_9388_) );
	NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf3), .B(_9344_), .C(_9388_), .Y(_9399_) );
	NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_8927_), .Y(_9410_) );
	NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_9410_), .B(_9267_), .Y(_9421_) );
	NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_9421_), .B(divider_divuResult_23_), .Y(_9432_) );
	NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_7709_), .B(_7731_), .C(_9147_), .Y(_9443_) );
	NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .B(_9432_), .C(_9443_), .Y(_9454_) );
	NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_9267_), .B(_9410_), .C(divider_divuResult_23_), .Y(_9465_) );
	OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_7929_), .B(_8280_), .C(_7709_), .Y(_9476_) );
	OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_9476_), .Y(_9487_) );
	NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf2), .B(_9487_), .C(_9465_), .Y(_9498_) );
	AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_9498_), .B(_9454_), .C(_9333_), .D(_9399_), .Y(_9509_) );
	AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .B(_9509_), .Y(_9520_) );
	OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .B(_8280_), .C(_8027_), .Y(_9531_) );
	INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(_9531_), .Y(_9542_) );
	OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_9542_), .Y(_9553_) );
	NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_8445_), .B(_8916_), .Y(_9564_) );
	NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_8379_), .C(_9564_), .Y(_9575_) );
	INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(_8445_), .Y(_9586_) );
	INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(_8643_), .Y(_9597_) );
	NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_8511_), .Y(_9608_) );
	AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_9597_), .B(_8522_), .C(_9608_), .Y(_9619_) );
	NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_8577_), .B(_8621_), .Y(_9630_) );
	OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_7478_), .Y(_9641_) );
	NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_8500_), .C(_9641_), .Y(_9652_) );
	OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_7380_), .C(_7467_), .Y(_9663_) );
	NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_8872_), .C(_9663_), .Y(_9674_) );
	NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_9652_), .B(_9674_), .Y(_9685_) );
	NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_8839_), .B(_9630_), .C(_9685_), .Y(_9696_) );
	AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_9696_), .B(_9619_), .C(_9586_), .Y(_9707_) );
	OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_8357_), .B(_9707_), .C(_8795_), .Y(_9718_) );
	NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_9575_), .B(_9718_), .Y(_9729_) );
	NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_8938_), .B(_8708_), .C(_9729_), .Y(_9740_) );
	AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_9740_), .B(_9553_), .C(_4100__bF_buf0), .Y(_9751_) );
	OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_9531_), .Y(_9762_) );
	OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_8357_), .B(_9707_), .C(_8379_), .Y(_9773_) );
	NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_8795_), .C(_9564_), .Y(_9784_) );
	NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_9784_), .B(_9773_), .Y(_9795_) );
	NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_8938_), .B(_8708_), .C(_9795_), .Y(_9806_) );
	AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_9806_), .B(_9762_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .Y(_9817_) );
	NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_9586_), .B(_8665_), .Y(_9828_) );
	NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_9564_), .B(_9828_), .Y(_9839_) );
	NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_9839_), .C(_8938_), .Y(_9850_) );
	OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_8346_), .Y(_9860_) );
	NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .B(_9850_), .C(_9860_), .Y(_9871_) );
	INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(_9839_), .Y(_9882_) );
	NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_8938_), .C(_9882_), .Y(_9893_) );
	OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_8773_), .Y(_9904_) );
	NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_9893_), .C(_9904_), .Y(_9915_) );
	NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_9871_), .B(_9915_), .Y(_9926_) );
	OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_9751_), .B(_9817_), .C(_9926_), .Y(_9937_) );
	OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_24_), .B(divider_divuResult_24_bF_buf3), .C(_8555_), .Y(_9948_) );
	OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .B(_9948_), .C(_8850_), .Y(_9959_) );
	XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_9959_), .B(_9685_), .Y(_9980_) );
	INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(_9980_), .Y(_9981_) );
	NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_9981_), .C(_8938_), .Y(_9992_) );
	OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_8883_), .B(divider_divuResult_23_), .C(_9992_), .Y(_10003_) );
	INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(_10003_), .Y(_10014_) );
	OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_8511_), .Y(_10025_) );
	NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf3), .B(_9992_), .C(_10025_), .Y(_10036_) );
	NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_8839_), .B(_9630_), .Y(_10047_) );
	NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_8632_), .B(_10047_), .Y(_10058_) );
	INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_10058_), .Y(_10069_) );
	NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_10069_), .C(_8938_), .Y(_10080_) );
	OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_9948_), .Y(_10091_) );
	NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_10080_), .C(_10091_), .Y(_10102_) );
	NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_10036_), .B(_10102_), .Y(_10113_) );
	OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_10014_), .C(_10113_), .Y(_10124_) );
	NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf7), .B(_9762_), .C(_9806_), .Y(_10135_) );
	INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(_10135_), .Y(_10146_) );
	OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_9147_), .B(_9729_), .C(_9762_), .Y(_10157_) );
	NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .B(_10157_), .Y(_10168_) );
	NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_9850_), .C(_9860_), .Y(_10179_) );
	INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(_10179_), .Y(_10190_) );
	AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_10190_), .B(_10168_), .C(_10146_), .Y(_10201_) );
	OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_10124_), .B(_9937_), .C(_10201_), .Y(_10212_) );
	NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_9037_), .B(_8960_), .Y(_10223_) );
	NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf2), .B(_9158_), .C(_9136_), .Y(_10234_) );
	NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .B(_9180_), .C(_9213_), .Y(_10245_) );
	NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_10245_), .B(_10234_), .C(_10223_), .Y(_10256_) );
	AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_9388_), .B(_9344_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .Y(_10267_) );
	NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_9245_), .B(_9322_), .Y(_10278_) );
	NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .B(_10278_), .Y(_10289_) );
	AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_9465_), .B(_9487_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .Y(_10300_) );
	OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_10300_), .B(_10267_), .C(_10289_), .Y(_10311_) );
	OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf4), .B(_8949_), .C(_8971__bF_buf5), .Y(_10322_) );
	INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(_10322_), .Y(_10333_) );
	AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_9213_), .B(_9180_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .Y(_10344_) );
	AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_10223_), .B(_10344_), .C(_10333_), .Y(_10355_) );
	OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_10256_), .B(_10311_), .C(_10355_), .Y(_10366_) );
	AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_9520_), .B(_10212_), .C(_10366_), .Y(_10377_) );
	NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .B(_9762_), .C(_9806_), .Y(_10388_) );
	NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf6), .B(_9553_), .C(_9740_), .Y(_10399_) );
	AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_9871_), .B(_9915_), .C(_10388_), .D(_10399_), .Y(_10410_) );
	XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf0), .B(divider_aOp_abs_23_), .Y(_10421_) );
	INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(_10421_), .Y(_10432_) );
	NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_10432_), .B(_8708_), .C(_8938_), .Y(_10441_) );
	OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_8533_), .Y(_10450_) );
	NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf6), .B(_10441_), .C(_10450_), .Y(_10460_) );
	AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_10450_), .B(_10441_), .C(_1768__bF_buf5), .Y(_10469_) );
	NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_22_), .B(_1746__bF_buf5), .Y(_10479_) );
	OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_10479_), .B(_10469_), .C(_10460_), .Y(_10487_) );
	NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .B(_9992_), .C(_10025_), .Y(_10497_) );
	OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_8883_), .Y(_10506_) );
	NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_9980_), .C(_8938_), .Y(_10516_) );
	NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_10516_), .C(_10506_), .Y(_10526_) );
	NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_10080_), .C(_10091_), .Y(_10535_) );
	OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_9015_), .C(_8894_), .Y(_10544_) );
	NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_8708_), .B(_10058_), .C(_8938_), .Y(_10554_) );
	NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_10554_), .C(_10544_), .Y(_10564_) );
	AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_10497_), .B(_10526_), .C(_10535_), .D(_10564_), .Y(_10574_) );
	NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_10574_), .B(_10487_), .C(_10410_), .Y(_10584_) );
	INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(_10584_), .Y(_10594_) );
	NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_10594_), .B(_9520_), .Y(_10604_) );
	AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_10377_), .B(_10604_), .C(_2185_), .Y(divider_divuResult_22_) );
	OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_7775_), .B(divider_divuResult_23_), .C(_2229__bF_buf1), .Y(_10623_) );
	INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .Y(_10633_) );
	NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_9509_), .B(_9234_), .Y(_10643_) );
	AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_10025_), .B(_9992_), .C(_2470__bF_buf0), .Y(_10653_) );
	OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_10102_), .B(_10653_), .C(_10036_), .Y(_10662_) );
	AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_9806_), .B(_9762_), .C(_4100__bF_buf5), .Y(_10663_) );
	OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_10179_), .B(_10663_), .C(_10135_), .Y(_10664_) );
	AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_10410_), .B(_10662_), .C(_10664_), .Y(_10665_) );
	NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf2), .B(_9245_), .C(_9322_), .Y(_10666_) );
	AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_9322_), .B(_9245_), .C(_4714__bF_buf1), .Y(_10667_) );
	OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_9147_), .B(_9421_), .C(_9487_), .Y(_10668_) );
	NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_10668_), .Y(_10669_) );
	AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_10666_), .B(_10669_), .C(_10667_), .Y(_10670_) );
	NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf4), .B(_10623_), .Y(_10671_) );
	OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_10671_), .B(_10234_), .C(_10322_), .Y(_10672_) );
	AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .B(_10670_), .C(_10672_), .Y(_10673_) );
	OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_10643_), .B(_10665_), .C(_10673_), .Y(_10674_) );
	NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_10584_), .B(_10643_), .Y(_10675_) );
	OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_10675_), .B(_10674_), .C(_10633_), .Y(_10676_) );
	AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_10676__bF_buf3), .B(_10623_), .C(_2240__bF_buf3), .Y(_10677_) );
	INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .Y(_10678_) );
	XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_10677_), .B(_10678__bF_buf5), .Y(_10679_) );
	NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_9224_), .B(_9169_), .Y(_10680_) );
	INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(_9509_), .Y(_10681_) );
	AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_10665_), .B(_10584_), .C(_10681_), .Y(_10682_) );
	OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_10670_), .B(_10682_), .C(_10680_), .Y(_10683_) );
	INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .Y(_1099_) );
	NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_10670_), .B(_10682_), .Y(_1100_) );
	NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1100_), .Y(_1101_) );
	NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_10683_), .B(divider_divuResult_22_), .C(_1101_), .Y(_1102_) );
	NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_9202_), .B(_9191_), .Y(_1103_) );
	OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_9147_), .B(_1103_), .C(_9180_), .Y(_1104_) );
	NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_10676__bF_buf2), .Y(_1105_) );
	AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1105_), .C(_8971__bF_buf3), .Y(_1106_) );
	INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(_10683_), .Y(_1107_) );
	NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .B(_10670_), .C(_10682_), .Y(_1108_) );
	OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_1107_), .C(divider_divuResult_22_), .Y(_1109_) );
	INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1110_) );
	NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .B(_10676__bF_buf1), .Y(_1111_) );
	AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1109_), .B(_1111_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .Y(_1112_) );
	OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1106_), .B(_1112_), .C(_10679_), .Y(_1113_) );
	NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_10278_), .B(_10676__bF_buf0), .Y(_1114_) );
	NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_9333_), .B(_9399_), .Y(_1115_) );
	INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .Y(_1116_) );
	NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_9454_), .B(_9498_), .Y(_1117_) );
	INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .Y(_1118_) );
	AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_10665_), .B(_10584_), .C(_1118_), .Y(_1119_) );
	OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_10300_), .B(_1119_), .C(_1116_), .Y(_1120_) );
	OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_10212_), .B(_10594_), .C(_1117_), .Y(_1121_) );
	NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_10669_), .C(_1121_), .Y(_1122_) );
	NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1120_), .B(_1122_), .C(divider_divuResult_22_), .Y(_1123_) );
	NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf1), .B(_1114_), .C(_1123_), .Y(_1124_) );
	OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_10300_), .B(_1119_), .C(_1115_), .Y(_1125_) );
	NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_10669_), .C(_1121_), .Y(_1126_) );
	NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .B(_1126_), .C(divider_divuResult_22_), .Y(_1127_) );
	INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(_10278_), .Y(_1128_) );
	NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_10676__bF_buf3), .Y(_1129_) );
	NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .B(_1129_), .C(_1127_), .Y(_1130_) );
	NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .B(_9509_), .C(_10212_), .Y(_1131_) );
	NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_10673_), .B(_1131_), .C(_10604_), .Y(_1132_) );
	NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_10584_), .C(_10665_), .Y(_1133_) );
	NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1121_), .Y(_1134_) );
	NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1132_), .C(_1134_), .Y(_1135_) );
	NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_9465_), .B(_9487_), .C(_10676__bF_buf2), .Y(_1136_) );
	NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_1135_), .C(_1136_), .Y(_1137_) );
	NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_10668_), .B(_10676__bF_buf1), .Y(_1138_) );
	INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .Y(_1139_) );
	NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1119_), .B(_1139_), .Y(_1140_) );
	NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1132_), .C(_1140_), .Y(_1141_) );
	NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf0), .B(_1138_), .C(_1141_), .Y(_1142_) );
	NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1142_), .Y(_1143_) );
	NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1124_), .B(_1130_), .C(_1143_), .Y(_1144_) );
	NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1113_), .Y(_1145_) );
	NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_10157_), .B(_10676__bF_buf0), .Y(_1146_) );
	NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_10388_), .B(_10399_), .Y(_1147_) );
	INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(_9926_), .Y(_1148_) );
	INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(_10653_), .Y(_1149_) );
	AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_10113_), .C(_10574_), .D(_10487_), .Y(_1150_) );
	OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1150_), .C(_10179_), .Y(_1151_) );
	NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1151_), .Y(_1152_) );
	INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .Y(_1153_) );
	NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_10421_), .B(_8719_), .C(_9015_), .Y(_1154_) );
	AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_8938_), .B(_8708_), .C(divider_aOp_abs_23_), .Y(_1155_) );
	NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .B(_1155_), .C(_1154_), .Y(_1156_) );
	OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1154_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .Y(_1157_) );
	INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_10479_), .Y(_1158_) );
	AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1158_), .C(_1156_), .Y(_1159_) );
	AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_10506_), .B(_10516_), .C(_2470__bF_buf7), .Y(_1160_) );
	AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_10025_), .B(_9992_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .Y(_1161_) );
	AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_10544_), .B(_10554_), .C(_2547__bF_buf2), .Y(_1162_) );
	AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_10091_), .B(_10080_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .Y(_1163_) );
	OAI22X1 OAI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1161_), .C(_1162_), .D(_1163_), .Y(_1164_) );
	OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_1159_), .C(_10124_), .Y(_1165_) );
	NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_9926_), .B(_1165_), .Y(_1166_) );
	NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_10179_), .C(_1166_), .Y(_1167_) );
	NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1152_), .B(_1167_), .Y(_1168_) );
	NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1132_), .C(_1168_), .Y(_1169_) );
	NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf0), .B(_1146_), .C(_1169_), .Y(_1170_) );
	NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_10179_), .C(_1166_), .Y(_1171_) );
	NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1151_), .Y(_1172_) );
	NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(_1171_), .Y(_1173_) );
	NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1132_), .C(_1173_), .Y(_1174_) );
	NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_9762_), .B(_9806_), .C(_10676__bF_buf3), .Y(_1175_) );
	NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_1175_), .C(_1174_), .Y(_1176_) );
	NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1150_), .Y(_1177_) );
	NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1166_), .Y(_1178_) );
	NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1178_), .C(_1132_), .Y(_1179_) );
	OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_8773_), .B(divider_divuResult_23_), .C(_9850_), .Y(_1180_) );
	NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(_10676__bF_buf2), .Y(_1181_) );
	NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(_1179_), .C(_1181_), .Y(_1182_) );
	INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .Y(_1183_) );
	NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1132_), .C(_1183_), .Y(_1184_) );
	NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_9850_), .B(_9860_), .C(_10676__bF_buf1), .Y(_1185_) );
	NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf4), .B(_1184_), .C(_1185_), .Y(_1186_) );
	NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1186_), .Y(_1187_) );
	NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_1176_), .C(_1187_), .Y(_1188_) );
	NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_10003_), .B(_10676__bF_buf0), .Y(_1189_) );
	NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_10497_), .B(_10526_), .Y(_1190_) );
	NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_1163_), .Y(_1191_) );
	OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(_1159_), .C(_10102_), .Y(_1192_) );
	XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1190_), .Y(_1193_) );
	NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1193_), .C(_1132_), .Y(_1194_) );
	NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_1194_), .C(_1189_), .Y(_1195_) );
	INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .Y(_1196_) );
	NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_10014_), .B(_10676__bF_buf3), .Y(_1197_) );
	INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .Y(_1198_) );
	XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1198_), .Y(_1199_) );
	NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1199_), .C(_1132_), .Y(_1200_) );
	NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .B(_1200_), .C(_1197_), .Y(_1201_) );
	OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_8894_), .B(divider_divuResult_23_), .C(_10080_), .Y(_1202_) );
	INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .Y(_1203_) );
	NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_10676__bF_buf2), .Y(_1204_) );
	XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_10487_), .B(_1191_), .Y(_1205_) );
	NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1205_), .C(_1132_), .Y(_1206_) );
	AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1206_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .Y(_1207_) );
	AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1201_), .C(_1196_), .Y(_1208_) );
	INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .Y(_1209_) );
	AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1184_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .Y(_1210_) );
	AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(_1176_), .C(_1209_), .Y(_1211_) );
	OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1188_), .C(_1211_), .Y(_1212_) );
	AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1129_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .Y(_1213_) );
	OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_10668_), .B(divider_divuResult_22_), .C(_1135_), .Y(_1214_) );
	NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .B(_1214_), .Y(_1215_) );
	AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_1130_), .C(_1213_), .Y(_1216_) );
	AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_2229__bF_buf0), .B(_9026_), .C(_10633_), .D(_1132_), .Y(_1217_) );
	OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf2), .B(_1217_), .C(_10678__bF_buf4), .Y(_1218_) );
	INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(_1218_), .Y(_1219_) );
	OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf1), .B(_8949_), .C(_10676__bF_buf1), .Y(_1220_) );
	NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .B(_2229__bF_buf4), .C(_1220_), .Y(_1221_) );
	AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1105_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .Y(_1222_) );
	AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_1221_), .C(_1219_), .Y(_1223_) );
	OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1216_), .B(_1113_), .C(_1223_), .Y(_1224_) );
	AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(_1212_), .C(_1224_), .Y(_1225_) );
	NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1154_), .Y(_1226_) );
	INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .Y(_1227_) );
	AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_10633_), .C(_1227_), .Y(_1228_) );
	NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_10469_), .B(_1156_), .Y(_1229_) );
	XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .B(_10479_), .Y(_1230_) );
	INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .Y(_1231_) );
	NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_10676__bF_buf0), .Y(_1232_) );
	OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1232_), .C(_2547__bF_buf1), .Y(_1233_) );
	OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1232_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .Y(_1234_) );
	NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_10676__bF_buf3), .Y(_1235_) );
	AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_10633_), .C(_1226_), .Y(_1236_) );
	OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1235_), .C(_2547__bF_buf0), .Y(_1237_) );
	NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1237_), .Y(_1238_) );
	INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_22_), .Y(_1239_) );
	NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .B(_1239_), .Y(_1240_) );
	INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1241_) );
	NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .B(_1241_), .Y(_1242_) );
	INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .Y(_1243_) );
	NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1243_), .C(_1132_), .Y(_1244_) );
	NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_10676__bF_buf2), .Y(_1245_) );
	NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_1244_), .C(_1245_), .Y(_1246_) );
	AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .B(_1244_), .C(_1768__bF_buf3), .Y(_1247_) );
	NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_21_), .B(_1746__bF_buf4), .Y(_1248_) );
	OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_1247_), .C(_1246_), .Y(_1249_) );
	NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1249_), .Y(_1250_) );
	AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1170_), .Y(_1251_) );
	NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .B(_1194_), .C(_1189_), .Y(_1252_) );
	NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf7), .B(_1200_), .C(_1197_), .Y(_1253_) );
	INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .Y(_1254_) );
	NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1254_), .C(_1132_), .Y(_1255_) );
	NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(_10676__bF_buf1), .Y(_1256_) );
	NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .B(_1255_), .C(_1256_), .Y(_1257_) );
	NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_1206_), .C(_1204_), .Y(_1258_) );
	AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1257_), .B(_1258_), .C(_1252_), .D(_1253_), .Y(_1259_) );
	NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1259_), .C(_1251_), .Y(_1260_) );
	AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1233_), .C(_1260_), .Y(_1261_) );
	NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(_1261_), .Y(_1262_) );
	AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_1262_), .C(_2503_), .Y(divider_divuResult_21_) );
	OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_10677_), .B(divider_divuResult_21_bF_buf4), .C(_2229__bF_buf3), .Y(_1263_) );
	NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .B(_1263_), .Y(_1264_) );
	INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .Y(_1265_) );
	INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .Y(_1266_) );
	NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1218_), .Y(_1267_) );
	NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .B(_1111_), .C(_1109_), .Y(_1268_) );
	NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf2), .B(_1105_), .C(_1102_), .Y(_1269_) );
	AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1269_), .C(_1267_), .Y(_1270_) );
	AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1114_), .C(_7204__bF_buf0), .Y(_1271_) );
	NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .B(_1271_), .Y(_1272_) );
	NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1143_), .C(_1270_), .Y(_1273_) );
	NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_1176_), .Y(_1274_) );
	AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1186_), .C(_1274_), .Y(_1275_) );
	OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(divider_divuResult_22_), .C(_1206_), .Y(_1276_) );
	NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf5), .B(_1276_), .Y(_1277_) );
	NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1201_), .Y(_1278_) );
	OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1277_), .B(_1278_), .C(_1195_), .Y(_1279_) );
	OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(divider_divuResult_22_), .C(_1184_), .Y(_1280_) );
	NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf3), .B(_1280_), .Y(_1281_) );
	OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1281_), .B(_1274_), .C(_1170_), .Y(_1282_) );
	AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1279_), .C(_1282_), .Y(_1283_) );
	OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_10676__bF_buf0), .B(_1134_), .C(_1138_), .Y(_1284_) );
	NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf6), .B(_1284_), .Y(_1285_) );
	OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1271_), .C(_1124_), .Y(_1286_) );
	OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .B(divider_divuResult_22_), .C(_1102_), .Y(_1287_) );
	NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf1), .B(_1287_), .Y(_1288_) );
	OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1288_), .C(_1218_), .Y(_1289_) );
	AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1270_), .C(_1289_), .Y(_1290_) );
	OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_1283_), .C(_1290_), .Y(_1291_) );
	INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .Y(_1292_) );
	AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .B(_1238_), .C(_1292_), .Y(_1293_) );
	NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1260_), .C(_1273_), .Y(_1294_) );
	OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1291_), .C(_1266_), .Y(_1295_) );
	OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf0), .B(_1217_), .C(_1295_), .Y(_1296_) );
	NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_2229__bF_buf2), .C(_1296_), .Y(_1297_) );
	NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1297_), .B(_1264_), .Y(_1298_) );
	NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1269_), .B(_1268_), .Y(_1299_) );
	INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .Y(_1300_) );
	INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .Y(_1301_) );
	OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1261_), .C(_1301_), .Y(_1302_) );
	AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1216_), .C(_1300_), .Y(_1303_) );
	AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_22_), .B(_1231_), .C(_1236_), .Y(_1304_) );
	NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_1304_), .Y(_1305_) );
	NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_1242_), .C(_1132_), .Y(_1306_) );
	NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_22_), .B(_10676__bF_buf3), .Y(_1307_) );
	AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1306_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .Y(_1308_) );
	NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .B(_1306_), .C(_1307_), .Y(_1309_) );
	INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .Y(_1310_) );
	AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1310_), .C(_1308_), .Y(_1311_) );
	OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .B(_1311_), .C(_1233_), .Y(_1312_) );
	NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1259_), .C(_1312_), .Y(_1313_) );
	AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .B(_1283_), .C(_1144_), .Y(_1314_) );
	NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1286_), .C(_1314_), .Y(_1315_) );
	OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1315_), .C(divider_divuResult_21_bF_buf3), .Y(_1316_) );
	INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .Y(_1317_) );
	NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1291_), .Y(_1318_) );
	OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1317_), .Y(_1319_) );
	NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf3), .B(_1319_), .C(_1316_), .Y(_1320_) );
	OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1314_), .C(_1299_), .Y(_1321_) );
	NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1216_), .C(_1302_), .Y(_1322_) );
	NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(divider_divuResult_21_bF_buf2), .C(_1321_), .Y(_1323_) );
	OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1287_), .Y(_1324_) );
	NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .B(_1324_), .C(_1323_), .Y(_1325_) );
	NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1325_), .C(_1298_), .Y(_1326_) );
	OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(divider_divuResult_22_), .C(_1123_), .Y(_1327_) );
	INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(_1327_), .Y(_1328_) );
	NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(divider_divuResult_21_bF_buf1), .Y(_1329_) );
	AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1142_), .C(_1283_), .D(_1313_), .Y(_1330_) );
	OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_1330_), .C(_1272_), .Y(_1331_) );
	INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1332_) );
	OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1212_), .B(_1261_), .C(_1143_), .Y(_1333_) );
	NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_1285_), .C(_1333_), .Y(_1334_) );
	AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .B(_1334_), .C(_1295_), .Y(_1335_) );
	OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1335_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .Y(_1336_) );
	OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1327_), .Y(_1337_) );
	NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1285_), .C(_1333_), .Y(_1338_) );
	OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_1330_), .C(_1332_), .Y(_1339_) );
	NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(divider_divuResult_21_bF_buf0), .C(_1339_), .Y(_1340_) );
	NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf0), .B(_1337_), .C(_1340_), .Y(_1341_) );
	INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1342_) );
	NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_1283_), .C(_1313_), .Y(_1343_) );
	NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1333_), .Y(_1344_) );
	NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(divider_divuResult_21_bF_buf4), .Y(_1345_) );
	OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(divider_divuResult_21_bF_buf3), .C(_1345_), .Y(_1346_) );
	OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .B(_1346_), .C(_1341_), .Y(_1347_) );
	NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1347_), .Y(_1348_) );
	NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf4), .B(_1263_), .Y(_1349_) );
	INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .Y(_1350_) );
	AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_1324_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .Y(_1351_) );
	AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1351_), .C(_1350_), .Y(_1352_) );
	OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(_1348_), .C(_1352_), .Y(_1353_) );
	NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .B(_1319_), .C(_1316_), .Y(_1354_) );
	NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf2), .B(_1324_), .C(_1323_), .Y(_1355_) );
	AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1297_), .C(_1355_), .D(_1354_), .Y(_1356_) );
	NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .B(_1337_), .C(_1340_), .Y(_1357_) );
	OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1335_), .C(_8971__bF_buf6), .Y(_1358_) );
	OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1214_), .Y(_1359_) );
	NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_1345_), .C(_1359_), .Y(_1360_) );
	AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1343_), .C(_1295_), .Y(_1361_) );
	NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(divider_divuResult_21_bF_buf2), .Y(_1362_) );
	OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1361_), .C(_7204__bF_buf5), .Y(_1363_) );
	AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1363_), .C(_1357_), .D(_1358_), .Y(_1364_) );
	AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1364_), .Y(_1365_) );
	OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_10676__bF_buf2), .B(_1173_), .C(_1146_), .Y(_1366_) );
	INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .Y(_1367_) );
	OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1367_), .Y(_1368_) );
	INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .Y(_1369_) );
	AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1259_), .C(_1279_), .Y(_1370_) );
	OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1370_), .C(_1281_), .Y(_1371_) );
	NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1251_), .B(_1371_), .Y(_1372_) );
	INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(_1259_), .Y(_1373_) );
	OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1293_), .C(_1208_), .Y(_1374_) );
	NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1374_), .Y(_1375_) );
	NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1281_), .C(_1375_), .Y(_1376_) );
	NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .B(divider_divuResult_21_bF_buf1), .C(_1372_), .Y(_1377_) );
	AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .B(_1368_), .C(_4714__bF_buf5), .Y(_1378_) );
	OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1366_), .Y(_1379_) );
	NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1251_), .B(_1281_), .C(_1375_), .Y(_1380_) );
	NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1371_), .Y(_1381_) );
	NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1380_), .B(divider_divuResult_21_bF_buf0), .C(_1381_), .Y(_1382_) );
	AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1379_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .Y(_1383_) );
	XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1187_), .Y(_1384_) );
	NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(divider_divuResult_21_bF_buf4), .Y(_1385_) );
	NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1295_), .Y(_1386_) );
	AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_1385_), .C(_4999__bF_buf6), .Y(_1387_) );
	NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1370_), .Y(_1388_) );
	NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1374_), .Y(_1389_) );
	OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1388_), .B(_1389_), .C(divider_divuResult_21_bF_buf3), .Y(_1390_) );
	INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .Y(_1391_) );
	NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1295_), .Y(_1392_) );
	AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1392_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .Y(_1393_) );
	OAI22X1 OAI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_1393_), .C(_1378_), .D(_1383_), .Y(_1394_) );
	INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(_1257_), .Y(_1395_) );
	INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .Y(_1396_) );
	NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_1396_), .Y(_1397_) );
	OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1293_), .C(_1277_), .Y(_1398_) );
	XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_1278_), .Y(_1399_) );
	OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_10014_), .B(divider_divuResult_22_), .C(_1194_), .Y(_1400_) );
	NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_1295_), .Y(_1401_) );
	OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1399_), .C(_1401_), .Y(_1402_) );
	NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .B(_1402_), .Y(_1403_) );
	OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1276_), .Y(_1404_) );
	XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1397_), .Y(_1405_) );
	NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(divider_divuResult_21_bF_buf2), .Y(_1406_) );
	AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1406_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .Y(_1407_) );
	INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .Y(_1408_) );
	NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1295_), .Y(_1409_) );
	NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_bF_buf1), .B(_1399_), .Y(_1410_) );
	AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(_1409_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .Y(_1411_) );
	OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_1407_), .C(_1403_), .Y(_1412_) );
	NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf4), .B(_1379_), .C(_1382_), .Y(_1413_) );
	INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .Y(_1414_) );
	NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_1368_), .C(_1377_), .Y(_1415_) );
	NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_1392_), .C(_1390_), .Y(_1416_) );
	INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .Y(_1417_) );
	AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_1417_), .C(_1414_), .Y(_1419_) );
	OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1394_), .C(_1419_), .Y(_1420_) );
	AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1365_), .B(_1420_), .C(_1353_), .Y(_1421_) );
	NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(_1379_), .C(_1382_), .Y(_1422_) );
	NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf3), .B(_1368_), .C(_1377_), .Y(_1423_) );
	NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .B(_1392_), .C(_1390_), .Y(_1424_) );
	NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_1385_), .C(_1386_), .Y(_1425_) );
	AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(_1425_), .C(_1422_), .D(_1423_), .Y(_1426_) );
	XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_1278_), .Y(_1427_) );
	NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_bF_buf0), .B(_1427_), .Y(_1428_) );
	NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_1401_), .C(_1428_), .Y(_1430_) );
	NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_1409_), .C(_1410_), .Y(_1431_) );
	INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .Y(_1432_) );
	NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(divider_divuResult_21_bF_buf4), .Y(_1433_) );
	INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .Y(_1434_) );
	OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_1318_), .C(_1434_), .Y(_1435_) );
	NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .B(_1433_), .C(_1435_), .Y(_1436_) );
	NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf6), .B(_1406_), .C(_1404_), .Y(_1437_) );
	AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(_1431_), .C(_1436_), .D(_1437_), .Y(_1438_) );
	AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1438_), .Y(_1439_) );
	NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1225_), .Y(_1441_) );
	OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1305_), .C(_1311_), .Y(_1442_) );
	NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1442_), .Y(_1443_) );
	NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1443_), .C(_1441_), .Y(_1444_) );
	OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1304_), .B(divider_divuResult_21_bF_buf3), .C(_1444_), .Y(_1445_) );
	NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .B(_1445_), .Y(_1446_) );
	OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_22_), .B(divider_divuResult_22_), .C(_1244_), .Y(_1447_) );
	INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .Y(_1448_) );
	NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1309_), .Y(_1449_) );
	XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .B(_1248_), .Y(_1450_) );
	NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1450_), .C(_1441_), .Y(_1452_) );
	OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(divider_divuResult_21_bF_buf2), .C(_1452_), .Y(_1453_) );
	OAI22X1 OAI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_1453_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .D(_1445_), .Y(_1454_) );
	NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1454_), .Y(_1455_) );
	INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .Y(_1456_) );
	NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1456_), .C(_1441_), .Y(_1457_) );
	NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_1304_), .B(_1295_), .Y(_1458_) );
	AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_1457_), .C(_2470__bF_buf4), .Y(_1459_) );
	NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1232_), .Y(_1460_) );
	NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_1295_), .Y(_1461_) );
	AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_1444_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .Y(_1463_) );
	INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .Y(_1464_) );
	NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(divider_divuResult_21_bF_buf1), .Y(_1465_) );
	NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(_1295_), .Y(_1466_) );
	AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1465_), .C(_2547__bF_buf6), .Y(_1467_) );
	NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1295_), .Y(_1468_) );
	AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1452_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .Y(_1469_) );
	OAI22X1 OAI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1463_), .C(_1467_), .D(_1469_), .Y(_1470_) );
	INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_21_), .Y(_1471_) );
	NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_1471_), .Y(_1472_) );
	OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_1472_), .C(divider_divuResult_21_bF_buf0), .Y(_1474_) );
	NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_21_), .B(_1295_), .Y(_1475_) );
	NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .B(_1475_), .C(_1474_), .Y(_1476_) );
	NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_20_), .B(_1746__bF_buf3), .Y(_1477_) );
	INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(_1477_), .Y(_1478_) );
	AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_1475_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .Y(_1479_) );
	OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1479_), .C(_1476_), .Y(_1480_) );
	OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1470_), .C(_1455_), .Y(_1481_) );
	NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1481_), .C(_1365_), .Y(_1482_) );
	AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1482_), .C(_3226_), .Y(divider_divuResult_20_) );
	INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .Y(_1484_) );
	AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1337_), .C(_8971__bF_buf5), .Y(_1485_) );
	NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf4), .B(_1345_), .C(_1359_), .Y(_1486_) );
	OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .B(_1485_), .C(_1341_), .Y(_1487_) );
	NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf3), .B(_1263_), .Y(_1488_) );
	OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1320_), .C(_1349_), .Y(_1489_) );
	AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1487_), .C(_1489_), .Y(_1490_) );
	NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_1356_), .Y(_1491_) );
	AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1428_), .B(_1401_), .C(_4100__bF_buf1), .Y(_1492_) );
	NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf5), .B(_1433_), .C(_1435_), .Y(_1493_) );
	NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf0), .B(_1401_), .C(_1428_), .Y(_1495_) );
	AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1495_), .C(_1492_), .Y(_1496_) );
	AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1379_), .C(_4714__bF_buf2), .Y(_1497_) );
	OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1497_), .C(_1413_), .Y(_1498_) );
	AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_1426_), .C(_1498_), .Y(_1499_) );
	OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1499_), .C(_1490_), .Y(_1500_) );
	NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1426_), .Y(_1501_) );
	NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_1444_), .C(_1461_), .Y(_1502_) );
	NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf3), .B(_1457_), .C(_1458_), .Y(_1503_) );
	NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_1452_), .C(_1468_), .Y(_1504_) );
	NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_1465_), .C(_1466_), .Y(_1506_) );
	AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1503_), .C(_1504_), .D(_1506_), .Y(_1507_) );
	NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_1472_), .Y(_1508_) );
	NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(divider_divuResult_21_bF_buf4), .Y(_1509_) );
	NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1295_), .Y(_1510_) );
	AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1510_), .B(_1509_), .C(_1768__bF_buf2), .Y(_1511_) );
	NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf1), .B(_1509_), .C(_1510_), .Y(_1512_) );
	AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1477_), .C(_1511_), .Y(_1513_) );
	AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1454_), .C(_1513_), .D(_1507_), .Y(_1514_) );
	NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1514_), .C(_1491_), .Y(_1515_) );
	OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1515_), .C(_3215_), .Y(_1517_) );
	AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf3), .B(_1263_), .C(_2240__bF_buf4), .Y(_1518_) );
	XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .B(_1484__bF_buf4), .Y(_1519_) );
	NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1355_), .B(_1354_), .Y(_1520_) );
	INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .Y(_1521_) );
	OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1514_), .C(_1499_), .Y(_1522_) );
	AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1364_), .C(_1487_), .Y(_1523_) );
	NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1523_), .Y(_1524_) );
	AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1521_), .Y(_1525_) );
	OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1525_), .C(divider_divuResult_20_bF_buf3), .Y(_1526_) );
	OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(divider_divuResult_21_bF_buf3), .C(_1323_), .Y(_1528_) );
	INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1529_) );
	AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1365_), .C(_1353_), .Y(_1530_) );
	OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1529_), .Y(_1531_) );
	NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf2), .B(_1531_), .C(_1526_), .Y(_1532_) );
	OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1521_), .Y(_1533_) );
	NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1523_), .Y(_1534_) );
	NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf2), .B(_1534_), .C(_1533_), .Y(_1535_) );
	OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1528_), .Y(_1536_) );
	NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .B(_1536_), .C(_1535_), .Y(_1537_) );
	NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(_1532_), .C(_1519_), .Y(_1539_) );
	OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(divider_divuResult_21_bF_buf2), .C(_1340_), .Y(_1540_) );
	OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1540_), .Y(_1541_) );
	NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1358_), .Y(_1542_) );
	NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1363_), .Y(_1543_) );
	NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .B(_1522_), .Y(_1544_) );
	NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .B(_1542_), .C(_1544_), .Y(_1545_) );
	INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .Y(_1546_) );
	INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .Y(_1547_) );
	NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1481_), .Y(_1548_) );
	AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1363_), .C(_1499_), .D(_1548_), .Y(_1550_) );
	OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .B(_1550_), .C(_1547_), .Y(_1551_) );
	NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf1), .B(_1545_), .C(_1551_), .Y(_1552_) );
	NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf1), .B(_1541_), .C(_1552_), .Y(_1553_) );
	INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .Y(_1554_) );
	OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .B(_1550_), .C(_1542_), .Y(_1555_) );
	NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .B(_1547_), .C(_1544_), .Y(_1556_) );
	AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1556_), .C(_1517__bF_buf2), .Y(_1557_) );
	OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_1557_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .Y(_1558_) );
	XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1543_), .Y(_1559_) );
	NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf0), .B(_1559_), .Y(_1561_) );
	OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1346_), .Y(_1562_) );
	NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .B(_1562_), .C(_1561_), .Y(_1563_) );
	XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1543_), .Y(_1564_) );
	NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf3), .B(_1564_), .Y(_1565_) );
	NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1359_), .C(_1517__bF_buf1), .Y(_1566_) );
	NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf4), .B(_1566_), .C(_1565_), .Y(_1567_) );
	NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_1567_), .Y(_1568_) );
	NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1568_), .C(_1558_), .Y(_1569_) );
	NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1539_), .Y(_1570_) );
	OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(divider_divuResult_21_bF_buf1), .C(_1382_), .Y(_1572_) );
	OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1572_), .Y(_1573_) );
	NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_1423_), .Y(_1574_) );
	NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1425_), .B(_1424_), .Y(_1575_) );
	INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .Y(_1576_) );
	OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .B(_1514_), .C(_1412_), .Y(_1577_) );
	NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1575_), .B(_1577_), .Y(_1578_) );
	NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_1416_), .C(_1578_), .Y(_1579_) );
	INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .Y(_1580_) );
	NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1578_), .Y(_1581_) );
	NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_1581_), .Y(_1583_) );
	NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf2), .B(_1579_), .C(_1583_), .Y(_1584_) );
	NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_1573_), .C(_1584_), .Y(_1585_) );
	INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .Y(_1586_) );
	OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1586_), .Y(_1587_) );
	OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .B(_1383_), .C(_1581_), .Y(_1588_) );
	NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_1416_), .C(_1578_), .Y(_1589_) );
	NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf1), .B(_1589_), .C(_1588_), .Y(_1590_) );
	NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_1587_), .C(_1590_), .Y(_1591_) );
	XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1575_), .Y(_1592_) );
	NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf0), .B(_1592_), .Y(_1594_) );
	NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1386_), .C(_1517__bF_buf0), .Y(_1595_) );
	NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .B(_1595_), .C(_1594_), .Y(_1596_) );
	OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1575_), .Y(_1597_) );
	NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1578_), .B(_1597_), .C(divider_divuResult_20_bF_buf3), .Y(_1598_) );
	OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(divider_divuResult_21_bF_buf0), .C(_1385_), .Y(_1599_) );
	OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1599_), .Y(_1600_) );
	NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf1), .B(_1600_), .C(_1598_), .Y(_1601_) );
	NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1596_), .B(_1601_), .Y(_1602_) );
	NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1591_), .C(_1602_), .Y(_1603_) );
	NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1403_), .Y(_1605_) );
	NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1437_), .Y(_1606_) );
	INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .Y(_1607_) );
	OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1607_), .B(_1514_), .C(_1493_), .Y(_1608_) );
	XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1605_), .Y(_1609_) );
	OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1402_), .Y(_1610_) );
	OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf3), .B(_1609_), .C(_1610_), .Y(_1611_) );
	NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_1611_), .Y(_1612_) );
	NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .B(_1611_), .Y(_1613_) );
	NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1435_), .C(_1517__bF_buf2), .Y(_1614_) );
	XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1607_), .Y(_1616_) );
	OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf1), .B(_1616_), .Y(_1617_) );
	AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_1614_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .Y(_1618_) );
	OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_1613_), .C(_1612_), .Y(_1619_) );
	AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1590_), .B(_1587_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .Y(_1620_) );
	AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .B(_1600_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .Y(_1621_) );
	AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1591_), .C(_1620_), .Y(_1622_) );
	OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(_1603_), .C(_1622_), .Y(_1623_) );
	NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .B(_1554_), .C(_1557_), .Y(_1624_) );
	AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1566_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .Y(_1625_) );
	AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1625_), .C(_1624_), .Y(_1627_) );
	NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .B(_1518_), .Y(_1628_) );
	AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_1536_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .Y(_1629_) );
	AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1519_), .C(_1628_), .Y(_1630_) );
	OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .B(_1627_), .C(_1630_), .Y(_1631_) );
	AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1623_), .C(_1631_), .Y(_1632_) );
	NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf3), .B(_1611_), .Y(_1633_) );
	AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_4999__bF_buf2), .Y(_1634_) );
	AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_1614_), .C(_4100__bF_buf7), .Y(_1635_) );
	OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf0), .B(_1616_), .C(_1614_), .Y(_1636_) );
	NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .B(_1636_), .Y(_1638_) );
	OAI22X1 OAI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(_1634_), .C(_1635_), .D(_1638_), .Y(_1639_) );
	NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .B(_1639_), .Y(_1640_) );
	NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1503_), .Y(_1641_) );
	OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_1469_), .C(_1513_), .Y(_1642_) );
	OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_1453_), .C(_1642_), .Y(_1643_) );
	OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1641_), .Y(_1644_) );
	OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1463_), .C(_1643_), .Y(_1645_) );
	NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .B(_1644_), .Y(_1646_) );
	MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_1646_), .S(_1517__bF_buf3), .Y(_1647_) );
	NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf4), .B(_1647_), .Y(_1649_) );
	INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .Y(_1650_) );
	AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf2), .B(_1445_), .Y(_1651_) );
	AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_1645_), .C(_1517__bF_buf1), .Y(_1652_) );
	OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1651_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .Y(_1653_) );
	INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(_1642_), .Y(_1654_) );
	NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_1506_), .Y(_1655_) );
	NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1513_), .Y(_1656_) );
	NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_1654_), .Y(_1657_) );
	OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1453_), .Y(_1658_) );
	OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf0), .B(_1657_), .C(_1658_), .Y(_1660_) );
	NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .B(_1660_), .Y(_1661_) );
	AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .B(_1653_), .C(_1650_), .Y(_1662_) );
	OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1654_), .B(_1656_), .C(divider_divuResult_20_bF_buf2), .Y(_1663_) );
	NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .B(_1658_), .C(_1663_), .Y(_1664_) );
	NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(divider_divuResult_20_bF_buf1), .Y(_1665_) );
	NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_1468_), .C(_1517__bF_buf3), .Y(_1666_) );
	NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_1666_), .C(_1665_), .Y(_1667_) );
	NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_1664_), .Y(_1668_) );
	NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(_1653_), .C(_1668_), .Y(_1669_) );
	NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1511_), .B(_1479_), .Y(_1671_) );
	XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(_1478_), .Y(_1672_) );
	INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .Y(_1673_) );
	OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_21_), .B(divider_divuResult_21_bF_buf4), .C(_1509_), .Y(_1674_) );
	OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1674_), .Y(_1675_) );
	OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf2), .B(_1673_), .C(_1675_), .Y(_1676_) );
	NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_1676_), .Y(_1677_) );
	INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_19_), .Y(_1678_) );
	INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_20_), .Y(_1679_) );
	NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(_1679_), .Y(_1680_) );
	NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1477_), .B(_1680_), .Y(_1682_) );
	NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1365_), .Y(_1683_) );
	NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1683_), .C(_1482_), .Y(_1684_) );
	NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_1682_), .C(_1684_), .Y(_1685_) );
	OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(_1679_), .Y(_1686_) );
	NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_1685_), .C(_1686_), .Y(_1687_) );
	OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_1530_), .C(divider_aOp_abs_20_), .Y(_1688_) );
	INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .Y(_1689_) );
	NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_1689_), .C(_1684_), .Y(_1690_) );
	NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf0), .B(_1690_), .C(_1688_), .Y(_1691_) );
	AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(_1678_), .C(_1687_), .D(_1691_), .Y(_1693_) );
	NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf7), .B(_1685_), .C(_1686_), .Y(_1694_) );
	OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_1676_), .C(_1694_), .Y(_1695_) );
	OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_1693_), .C(_1677_), .Y(_1696_) );
	OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .B(_1696_), .C(_1662_), .Y(_1697_) );
	NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1640_), .B(_1570_), .C(_1697_), .Y(_1698_) );
	AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1698_), .C(_8697__bF_buf2), .Y(divider_divuResult_19_) );
	INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(_2174_), .Y(_1699_) );
	NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .B(divider_divuResult_19_bF_buf5), .Y(_1700_) );
	OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf3), .B(_1700_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .Y(_1701_) );
	INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(_1518_), .Y(_1703_) );
	AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1698_), .Y(_1704_) );
	OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf1), .B(_1704__bF_buf3), .C(_1703_), .Y(_1705_) );
	NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf3), .B(_2229__bF_buf1), .C(_1705_), .Y(_1706_) );
	NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1706_), .B(_1701_), .Y(_1707_) );
	OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(divider_divuResult_20_bF_buf0), .C(_1535_), .Y(_1708_) );
	NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .B(_1708_), .Y(_1709_) );
	NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf1), .B(_1536_), .C(_1535_), .Y(_1710_) );
	NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1710_), .B(_1709_), .Y(_1711_) );
	INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .Y(_1712_) );
	INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .Y(_1714_) );
	AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_1591_), .B(_1585_), .Y(_1715_) );
	NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf3), .B(_1609_), .Y(_1716_) );
	OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(divider_divuResult_20_bF_buf2), .C(_1716_), .Y(_1717_) );
	NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .B(_1717_), .Y(_1718_) );
	NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_1611_), .Y(_1719_) );
	NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .B(_1636_), .Y(_1720_) );
	NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf6), .B(_1614_), .C(_1617_), .Y(_1721_) );
	AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1720_), .B(_1721_), .C(_1719_), .D(_1718_), .Y(_1722_) );
	NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1722_), .C(_1715_), .Y(_1723_) );
	NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_1647_), .Y(_1725_) );
	OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1651_), .C(_1735__bF_buf3), .Y(_1726_) );
	AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .B(_1667_), .C(_1726_), .D(_1725_), .Y(_1727_) );
	NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .B(_1690_), .C(_1688_), .Y(_1728_) );
	NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_19_), .B(_1746__bF_buf2), .Y(_1729_) );
	INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .Y(_1730_) );
	NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1694_), .C(_1728_), .Y(_1731_) );
	MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1672_), .S(_1517__bF_buf1), .Y(_1732_) );
	OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_1679_), .B(divider_divuResult_20_bF_buf1), .C(_1690_), .Y(_1733_) );
	AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1768__bF_buf6), .C(_2547__bF_buf4), .D(_1732_), .Y(_1734_) );
	AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .B(_1676_), .C(_1731_), .D(_1734_), .Y(_1736_) );
	NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1736_), .Y(_1737_) );
	AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1662_), .C(_1723_), .Y(_1738_) );
	OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1738_), .C(_1714_), .Y(_1739_) );
	AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1627_), .C(_1712_), .Y(_1740_) );
	AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1640_), .C(_1623_), .Y(_1741_) );
	OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1741_), .C(_1627_), .Y(_1742_) );
	NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1742_), .Y(_1743_) );
	OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_1743_), .C(divider_divuResult_19_bF_buf4), .Y(_1744_) );
	OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf3), .B(_1708_), .Y(_1745_) );
	NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf3), .B(_1745_), .C(_1744_), .Y(_1747_) );
	NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1742_), .Y(_1748_) );
	NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1712_), .B(_1627_), .C(_1739_), .Y(_1749_) );
	NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf2), .B(_1749_), .C(_1748_), .Y(_1750_) );
	OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf0), .B(_1704__bF_buf2), .C(_1708_), .Y(_1751_) );
	NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .B(_1751_), .C(_1750_), .Y(_1752_) );
	NAND3X1 NAND3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1707_), .C(_1747_), .Y(_1753_) );
	AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1552_), .C(divider_divuResult_19_bF_buf1), .Y(_1754_) );
	INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf0), .Y(_1755_) );
	NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1558_), .Y(_1756_) );
	INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .Y(_1758_) );
	INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .Y(_1759_) );
	NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1640_), .B(_1697_), .Y(_1760_) );
	AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_1567_), .C(_1759_), .D(_1760_), .Y(_1761_) );
	OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1761_), .C(_1758_), .Y(_1762_) );
	INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .Y(_1763_) );
	OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1738_), .C(_1568_), .Y(_1764_) );
	NAND3X1 NAND3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .B(_1763_), .C(_1764_), .Y(_1765_) );
	AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1762_), .B(_1765_), .C(_1755_), .Y(_1766_) );
	NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .B(_1754_), .C(_1766_), .Y(_1767_) );
	OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf0), .B(_1559_), .C(_1566_), .Y(_1769_) );
	INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .Y(_1770_) );
	AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(_1770_), .Y(_1771_) );
	OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(_1771_), .C(divider_divuResult_19_bF_buf5), .Y(_1772_) );
	OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(divider_divuResult_19_bF_buf4), .C(_1772_), .Y(_1773_) );
	NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .B(_1773_), .Y(_1774_) );
	OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .B(_1766_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .Y(_1775_) );
	AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1775_), .B(_1774_), .C(_1767_), .Y(_1776_) );
	NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf2), .B(_1700_), .Y(_1777_) );
	NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .B(_1777_), .Y(_1778_) );
	AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1750_), .B(_1751_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .Y(_1780_) );
	AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1707_), .C(_1778_), .Y(_1781_) );
	OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1776_), .C(_1781_), .Y(_1782_) );
	INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .Y(_1783_) );
	NAND3X1 NAND3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1763_), .C(_1764_), .Y(_1784_) );
	OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1761_), .C(_1756_), .Y(_1785_) );
	NAND3X1 NAND3X1_376 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf3), .B(_1784_), .C(_1785_), .Y(_1786_) );
	NAND3X1 NAND3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf0), .B(_1783_), .C(_1786_), .Y(_1787_) );
	INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1788_) );
	OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf3), .B(_1704__bF_buf1), .C(_1788_), .Y(_1789_) );
	NAND3X1 NAND3X1_378 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .B(_1789_), .C(_1772_), .Y(_1791_) );
	NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1770_), .B(_1741_), .Y(_1792_) );
	NAND3X1 NAND3X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1764_), .B(_1792_), .C(divider_divuResult_19_bF_buf2), .Y(_1793_) );
	OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf2), .B(_1704__bF_buf0), .C(_1769_), .Y(_1794_) );
	NAND3X1 NAND3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf0), .B(_1793_), .C(_1794_), .Y(_1795_) );
	NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1795_), .B(_1791_), .Y(_1796_) );
	NAND3X1 NAND3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1787_), .B(_1796_), .C(_1775_), .Y(_1797_) );
	NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_1753_), .Y(_1798_) );
	INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .Y(_1799_) );
	INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .Y(_1800_) );
	AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1722_), .C(_1800_), .Y(_1802_) );
	NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1802_), .Y(_1803_) );
	OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1803_), .C(_1715_), .Y(_1804_) );
	NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1591_), .Y(_1805_) );
	INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_1806_) );
	INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .Y(_1807_) );
	NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_1807_), .Y(_1808_) );
	NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1649_), .Y(_1809_) );
	OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .B(_1809_), .C(_1649_), .Y(_1810_) );
	AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1727_), .C(_1810_), .Y(_1811_) );
	OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1811_), .C(_1619_), .Y(_1813_) );
	NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1813_), .Y(_1814_) );
	NAND3X1 NAND3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(_1806_), .C(_1814_), .Y(_1815_) );
	NAND3X1 NAND3X1_383 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf1), .B(_1815_), .C(_1804_), .Y(_1816_) );
	OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_1586_), .B(divider_divuResult_20_bF_buf0), .C(_1584_), .Y(_1817_) );
	INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(_1817_), .Y(_1818_) );
	OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf1), .B(_1704__bF_buf3), .C(_1818_), .Y(_1819_) );
	NAND3X1 NAND3X1_384 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_1819_), .C(_1816_), .Y(_1820_) );
	AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1816_), .B(_1819_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .Y(_1821_) );
	OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1517__bF_buf3), .B(_1592_), .C(_1600_), .Y(_1822_) );
	AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_1799_), .Y(_1824_) );
	OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_1824_), .C(divider_divuResult_19_bF_buf0), .Y(_1825_) );
	OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_1822_), .B(divider_divuResult_19_bF_buf5), .C(_1825_), .Y(_1826_) );
	NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .B(_1826_), .Y(_1827_) );
	OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1821_), .C(_1820_), .Y(_1828_) );
	OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf0), .B(_1704__bF_buf2), .C(_1817_), .Y(_1829_) );
	NAND3X1 NAND3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(_1806_), .C(_1814_), .Y(_1830_) );
	OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1803_), .C(_1805_), .Y(_1831_) );
	NAND3X1 NAND3X1_386 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf4), .B(_1830_), .C(_1831_), .Y(_1832_) );
	NAND3X1 NAND3X1_387 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf3), .B(_1829_), .C(_1832_), .Y(_1833_) );
	INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(_1822_), .Y(_1835_) );
	OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf3), .B(_1704__bF_buf1), .C(_1835_), .Y(_1836_) );
	NAND3X1 NAND3X1_388 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .B(_1836_), .C(_1825_), .Y(_1837_) );
	OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf2), .B(_1704__bF_buf0), .C(_1822_), .Y(_1838_) );
	NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_1802_), .Y(_1839_) );
	NAND3X1 NAND3X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1814_), .C(divider_divuResult_19_bF_buf3), .Y(_1840_) );
	NAND3X1 NAND3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf2), .B(_1840_), .C(_1838_), .Y(_1841_) );
	NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .B(_1837_), .Y(_1842_) );
	NAND3X1 NAND3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_1820_), .C(_1833_), .Y(_1843_) );
	OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf1), .B(_1704__bF_buf3), .C(_1717_), .Y(_1844_) );
	NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_1718_), .Y(_1846_) );
	INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(_1846_), .Y(_1847_) );
	INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .Y(_1848_) );
	OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_1638_), .C(_1697_), .Y(_1849_) );
	OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(_1848_), .C(_1849_), .Y(_1850_) );
	NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1847_), .B(_1850_), .Y(_1851_) );
	INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .Y(_1852_) );
	AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_1852_), .C(_1846_), .Y(_1853_) );
	OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_1851_), .C(divider_divuResult_19_bF_buf2), .Y(_1854_) );
	NAND3X1 NAND3X1_392 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_1844_), .C(_1854_), .Y(_1855_) );
	AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1854_), .B(_1844_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .Y(_1857_) );
	NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(_1720_), .Y(_1858_) );
	AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1858_), .Y(_1859_) );
	NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1858_), .B(_1697_), .Y(_1860_) );
	OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_1859_), .B(_1860_), .C(divider_divuResult_19_bF_buf1), .Y(_1861_) );
	OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(divider_divuResult_19_bF_buf0), .C(_1861_), .Y(_1862_) );
	NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .B(_1862_), .Y(_1863_) );
	OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_1857_), .C(_1855_), .Y(_1864_) );
	OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1843_), .C(_1828_), .Y(_1865_) );
	AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1865_), .C(_1782_), .Y(_1866_) );
	AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1854_), .B(_1844_), .C(_4714__bF_buf0), .Y(_1868_) );
	OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf0), .B(_1704__bF_buf2), .C(_1611_), .Y(_1869_) );
	AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_1852_), .C(_1847_), .Y(_1870_) );
	NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1846_), .B(_1850_), .Y(_1871_) );
	OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_1870_), .B(_1871_), .C(divider_divuResult_19_bF_buf5), .Y(_1872_) );
	AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(_1869_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .Y(_1873_) );
	NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf0), .B(_1862_), .Y(_1874_) );
	NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_1859_), .Y(_1875_) );
	NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(divider_divuResult_19_bF_buf4), .Y(_1876_) );
	OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(divider_divuResult_19_bF_buf3), .C(_1876_), .Y(_1877_) );
	NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_1877_), .Y(_1879_) );
	OAI22X1 OAI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .B(_1874_), .C(_1868_), .D(_1873_), .Y(_1880_) );
	NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1880_), .B(_1843_), .Y(_1881_) );
	NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_1732_), .Y(_1882_) );
	NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1677_), .B(_1882_), .Y(_1883_) );
	INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .Y(_1884_) );
	OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .B(_1884_), .C(_1731_), .Y(_1885_) );
	XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_1883_), .Y(_1886_) );
	NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(divider_divuResult_19_bF_buf2), .Y(_1887_) );
	OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf3), .B(_1704__bF_buf1), .C(_1676_), .Y(_1888_) );
	NAND3X1 NAND3X1_393 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_1887_), .C(_1888_), .Y(_1890_) );
	OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf2), .B(_1704__bF_buf0), .C(_1732_), .Y(_1891_) );
	INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .Y(_1892_) );
	NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(divider_divuResult_19_bF_buf1), .Y(_1893_) );
	NAND3X1 NAND3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_1893_), .C(_1891_), .Y(_1894_) );
	NAND3X1 NAND3X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(_1687_), .C(_1691_), .Y(_1895_) );
	AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_1895_), .B(_1731_), .Y(_1896_) );
	INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .Y(_1897_) );
	NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(divider_divuResult_19_bF_buf0), .Y(_1898_) );
	OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf1), .B(_1704__bF_buf3), .C(_1884_), .Y(_1899_) );
	NAND3X1 NAND3X1_396 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_1898_), .C(_1899_), .Y(_1901_) );
	OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf0), .B(_1704__bF_buf2), .C(_1733_), .Y(_1902_) );
	NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(divider_divuResult_19_bF_buf5), .Y(_1903_) );
	NAND3X1 NAND3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_1903_), .C(_1902_), .Y(_1904_) );
	AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .B(_1894_), .C(_1901_), .D(_1904_), .Y(_1905_) );
	NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf1), .B(_1678_), .Y(_1906_) );
	NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(divider_aOp_abs_19_), .Y(_1907_) );
	OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(_1907_), .C(divider_divuResult_19_bF_buf4), .Y(_1908_) );
	OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf3), .B(_1704__bF_buf1), .C(_1678_), .Y(_1909_) );
	NAND3X1 NAND3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_1908_), .C(_1909_), .Y(_1910_) );
	AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1909_), .B(_1908_), .C(_1768__bF_buf4), .Y(_1911_) );
	NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_18_), .B(_1746__bF_buf0), .Y(_1912_) );
	OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_1911_), .C(_1910_), .Y(_1913_) );
	NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_1913_), .Y(_1914_) );
	INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .Y(_1915_) );
	OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf2), .B(_1704__bF_buf0), .C(_1915_), .Y(_1916_) );
	AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1668_), .C(_1661_), .Y(_1917_) );
	XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1917_), .B(_1809_), .Y(_1918_) );
	NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(divider_divuResult_19_bF_buf3), .Y(_1919_) );
	NAND3X1 NAND3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf5), .B(_1919_), .C(_1916_), .Y(_1920_) );
	OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_1732_), .B(divider_divuResult_19_bF_buf2), .C(_1887_), .Y(_1923_) );
	NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .B(_1923_), .Y(_1924_) );
	AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1919_), .C(_4100__bF_buf4), .Y(_1925_) );
	XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1668_), .Y(_1926_) );
	INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .Y(_1927_) );
	NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_1927_), .B(divider_divuResult_19_bF_buf1), .Y(_1928_) );
	OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf1), .B(_1704__bF_buf3), .C(_1660_), .Y(_1929_) );
	NAND3X1 NAND3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_1928_), .C(_1929_), .Y(_1930_) );
	OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1925_), .C(_1920_), .Y(_1931_) );
	OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(divider_divuResult_19_bF_buf0), .C(_1898_), .Y(_1932_) );
	OAI22X1 OAI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_1932_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .D(_1923_), .Y(_1934_) );
	AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_1934_), .C(_1931_), .Y(_1935_) );
	OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(divider_divuResult_19_bF_buf5), .C(_1919_), .Y(_1936_) );
	NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .B(_1936_), .Y(_1937_) );
	NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(divider_divuResult_19_bF_buf4), .Y(_1938_) );
	OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(divider_divuResult_19_bF_buf3), .C(_1938_), .Y(_1939_) );
	OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_1939_), .C(_1937_), .Y(_1940_) );
	AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_1940_), .C(_1914_), .D(_1935_), .Y(_1941_) );
	NAND3X1 NAND3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1881_), .C(_1941_), .Y(_1942_) );
	AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(_1866_), .C(_1699__bF_buf4), .Y(divider_divuResult_18_) );
	INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .Y(_1944_) );
	NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1757__bF_buf1), .Y(_1945_) );
	INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .Y(_1946_) );
	OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(divider_divuResult_18_bF_buf5), .C(_2229__bF_buf0), .Y(_1947_) );
	INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .Y(_1948_) );
	XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .Y(_1949_) );
	NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(_1748_), .Y(_1950_) );
	OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1950_), .C(_1751_), .Y(_1951_) );
	NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .B(_1951_), .Y(_1952_) );
	INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(_1951_), .Y(_1953_) );
	NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf2), .B(_1953_), .Y(_1955_) );
	INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .Y(_1956_) );
	INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .Y(_1957_) );
	OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(_1880_), .Y(_1958_) );
	AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_1913_), .B(_1905_), .Y(_1959_) );
	NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .B(_1936_), .Y(_1960_) );
	OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_8697__bF_buf0), .B(_1704__bF_buf2), .C(_1807_), .Y(_1961_) );
	AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .B(_1938_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .Y(_1962_) );
	AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(_1937_), .C(_1960_), .Y(_1963_) );
	AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_1893_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .Y(_1964_) );
	AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .B(_1903_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .Y(_1966_) );
	OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_1966_), .C(_1924_), .Y(_1967_) );
	NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_1963_), .Y(_1968_) );
	OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .B(_1936_), .C(_1940_), .Y(_1969_) );
	OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_1968_), .B(_1959_), .C(_1969_), .Y(_1970_) );
	OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(_1970_), .C(_1957_), .Y(_1971_) );
	NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1971_), .Y(_1972_) );
	AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(_1955_), .C(_1776_), .D(_1972_), .Y(_1973_) );
	NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1747_), .Y(_1974_) );
	INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .Y(_1975_) );
	INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(_1776_), .Y(_1977_) );
	NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_1914_), .B(_1935_), .Y(_1978_) );
	NAND3X1 NAND3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1881_), .C(_1978_), .Y(_1979_) );
	AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1979_), .B(_1957_), .C(_1797_), .Y(_1980_) );
	NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1975_), .B(_1977_), .C(_1980_), .Y(_1981_) );
	OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_1981_), .B(_1973_), .C(divider_divuResult_18_bF_buf4), .Y(_1982_) );
	AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(_1866_), .Y(_1983_) );
	OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf3), .B(_1983__bF_buf4), .C(_1953_), .Y(_1984_) );
	NAND3X1 NAND3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf2), .B(_1984_), .C(_1982_), .Y(_1985_) );
	OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_1977_), .B(_1980_), .C(_1975_), .Y(_1986_) );
	NAND3X1 NAND3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .B(_1776_), .C(_1972_), .Y(_1988_) );
	NAND3X1 NAND3X1_405 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf3), .B(_1986_), .C(_1988_), .Y(_1989_) );
	OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf2), .B(_1983__bF_buf3), .C(_1951_), .Y(_1990_) );
	NAND3X1 NAND3X1_406 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .B(_1990_), .C(_1989_), .Y(_1991_) );
	NAND3X1 NAND3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .B(_1991_), .C(_1985_), .Y(_1992_) );
	NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1787_), .B(_1775_), .Y(_1993_) );
	INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .Y(_1994_) );
	INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(_1796_), .Y(_1995_) );
	AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1979_), .B(_1957_), .C(_1995_), .Y(_1996_) );
	OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_1996_), .C(_1994_), .Y(_1997_) );
	INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .Y(_1999_) );
	NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1796_), .B(_1971_), .Y(_2000_) );
	NAND3X1 NAND3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(_1993_), .C(_2000_), .Y(_2001_) );
	NAND3X1 NAND3X1_409 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf2), .B(_1997_), .C(_2001_), .Y(_2002_) );
	NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .B(_1766_), .Y(_2003_) );
	OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf1), .B(_1983__bF_buf2), .C(_2003_), .Y(_2004_) );
	AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2004_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .Y(_2005_) );
	NAND3X1 NAND3X1_410 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .B(_2004_), .C(_2002_), .Y(_2006_) );
	NAND3X1 NAND3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .B(_1957_), .C(_1979_), .Y(_2007_) );
	NAND3X1 NAND3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .B(_2000_), .C(divider_divuResult_18_bF_buf1), .Y(_2008_) );
	INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(_1773_), .Y(_2010_) );
	OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf0), .B(_1983__bF_buf1), .C(_2010_), .Y(_2011_) );
	AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2011_), .B(_2008_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .Y(_2012_) );
	AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_2012_), .C(_2005_), .Y(_2013_) );
	NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf2), .B(_1948_), .Y(_2014_) );
	AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1989_), .B(_1990_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .Y(_2015_) );
	AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_2015_), .B(_1949_), .C(_2014_), .Y(_2016_) );
	OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2013_), .B(_1992_), .C(_2016_), .Y(_2017_) );
	INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(_2003_), .Y(_2018_) );
	OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf4), .B(_1983__bF_buf0), .C(_2018_), .Y(_2019_) );
	OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_1996_), .C(_1993_), .Y(_2021_) );
	NAND3X1 NAND3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(_1994_), .C(_2000_), .Y(_2022_) );
	NAND3X1 NAND3X1_414 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf0), .B(_2021_), .C(_2022_), .Y(_2023_) );
	NAND3X1 NAND3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf1), .B(_2019_), .C(_2023_), .Y(_2024_) );
	INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .Y(_2025_) );
	OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_2025_), .C(divider_divuResult_18_bF_buf5), .Y(_2026_) );
	OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf3), .B(_1983__bF_buf4), .C(_1773_), .Y(_2027_) );
	NAND3X1 NAND3X1_416 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .B(_2027_), .C(_2026_), .Y(_2028_) );
	NAND3X1 NAND3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_2008_), .C(_2011_), .Y(_2029_) );
	NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2029_), .B(_2028_), .Y(_2030_) );
	NAND3X1 NAND3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2006_), .C(_2030_), .Y(_2032_) );
	NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_1992_), .Y(_2033_) );
	OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(divider_divuResult_19_bF_buf2), .C(_1832_), .Y(_2034_) );
	OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf2), .B(_1983__bF_buf3), .C(_2034_), .Y(_2035_) );
	INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .Y(_2036_) );
	NAND3X1 NAND3X1_419 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .B(_1829_), .C(_1832_), .Y(_2037_) );
	NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf2), .B(_2034_), .Y(_2038_) );
	NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2038_), .Y(_2039_) );
	OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_1880_), .B(_1970_), .C(_1864_), .Y(_2040_) );
	NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_2040_), .Y(_2041_) );
	NAND3X1 NAND3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_2039_), .C(_2041_), .Y(_2043_) );
	INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .Y(_2044_) );
	INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .Y(_2045_) );
	INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(_1880_), .Y(_2046_) );
	NAND3X1 NAND3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(_1969_), .C(_1978_), .Y(_2047_) );
	AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2047_), .B(_1864_), .C(_2045_), .Y(_2048_) );
	OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_2048_), .C(_2044_), .Y(_2049_) );
	NAND3X1 NAND3X1_422 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf4), .B(_2049_), .C(_2043_), .Y(_2050_) );
	NAND3X1 NAND3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf5), .B(_2035_), .C(_2050_), .Y(_2051_) );
	INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .Y(_2052_) );
	OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf1), .B(_1983__bF_buf2), .C(_2052_), .Y(_2054_) );
	OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_2048_), .C(_2039_), .Y(_2055_) );
	NAND3X1 NAND3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_2044_), .C(_2041_), .Y(_2056_) );
	NAND3X1 NAND3X1_425 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf3), .B(_2055_), .C(_2056_), .Y(_2057_) );
	NAND3X1 NAND3X1_426 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .B(_2054_), .C(_2057_), .Y(_2058_) );
	OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(divider_divuResult_19_bF_buf1), .C(_1872_), .Y(_2059_) );
	NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf6), .B(_1877_), .Y(_2060_) );
	OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_2059_), .C(_2060_), .Y(_2061_) );
	AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_2061_), .C(_2046_), .D(_1941_), .Y(_2062_) );
	AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_2045_), .Y(_2063_) );
	OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(_2063_), .C(divider_divuResult_18_bF_buf2), .Y(_2065_) );
	OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf0), .B(_1983__bF_buf1), .C(_1826_), .Y(_2066_) );
	NAND3X1 NAND3X1_427 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .B(_2066_), .C(_2065_), .Y(_2067_) );
	NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2062_), .Y(_2068_) );
	NAND3X1 NAND3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_2041_), .C(divider_divuResult_18_bF_buf1), .Y(_2069_) );
	INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .Y(_2070_) );
	OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf4), .B(_1983__bF_buf0), .C(_2070_), .Y(_2071_) );
	NAND3X1 NAND3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf1), .B(_2069_), .C(_2071_), .Y(_2072_) );
	NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2072_), .B(_2067_), .Y(_2073_) );
	NAND3X1 NAND3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2051_), .B(_2058_), .C(_2073_), .Y(_2074_) );
	OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(divider_divuResult_19_bF_buf0), .C(_1854_), .Y(_2076_) );
	INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .Y(_2077_) );
	INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(_1873_), .Y(_2078_) );
	NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_2077_), .B(_2078_), .Y(_2079_) );
	INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(_2079_), .Y(_2080_) );
	NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .B(_1874_), .Y(_2081_) );
	OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .B(_1970_), .C(_2060_), .Y(_2082_) );
	OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_2082_), .B(_2080_), .Y(_2083_) );
	NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .B(_1970_), .Y(_2084_) );
	OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_2084_), .C(_2080_), .Y(_2085_) );
	NAND3X1 NAND3X1_431 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf0), .B(_2085_), .C(_2083_), .Y(_2087_) );
	OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2076_), .B(divider_divuResult_18_bF_buf5), .C(_2087_), .Y(_2088_) );
	NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .B(_2088_), .Y(_2089_) );
	OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf3), .B(_1983__bF_buf4), .C(_2076_), .Y(_2090_) );
	OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .B(_1873_), .C(_2082_), .Y(_2091_) );
	OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_2082_), .B(_2079_), .Y(_2092_) );
	NAND3X1 NAND3X1_432 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf4), .B(_2091_), .C(_2092_), .Y(_2093_) );
	AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_2090_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .Y(_2094_) );
	OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf2), .B(_1983__bF_buf3), .C(_1877_), .Y(_2095_) );
	AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_1970_), .B(_2081_), .Y(_2096_) );
	NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2096_), .Y(_2098_) );
	NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf3), .B(_2098_), .Y(_2099_) );
	AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2095_), .B(_2099_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .Y(_2100_) );
	OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .B(_2094_), .C(_2089_), .Y(_2101_) );
	AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(_2054_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .Y(_2102_) );
	AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_2069_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .Y(_2103_) );
	AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(_2103_), .C(_2102_), .Y(_2104_) );
	OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .B(_2074_), .C(_2104_), .Y(_2105_) );
	AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2033_), .C(_2017_), .Y(_2106_) );
	AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_2090_), .C(_7204__bF_buf1), .Y(_2107_) );
	OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf1), .B(_1983__bF_buf2), .C(_2059_), .Y(_2109_) );
	AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(_2109_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .Y(_2110_) );
	AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2095_), .B(_2099_), .C(_4714__bF_buf6), .Y(_2111_) );
	OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2096_), .C(divider_divuResult_18_bF_buf2), .Y(_2112_) );
	OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf0), .B(_1983__bF_buf1), .C(_1862_), .Y(_2113_) );
	AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2112_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .Y(_2114_) );
	OAI22X1 OAI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2114_), .C(_2107_), .D(_2110_), .Y(_2115_) );
	NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(_2074_), .Y(_2116_) );
	OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf4), .B(_1983__bF_buf0), .C(_1936_), .Y(_2117_) );
	NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .B(_1960_), .Y(_2118_) );
	INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(_1939_), .Y(_2120_) );
	NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .B(_2120_), .Y(_2121_) );
	NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_2121_), .Y(_2122_) );
	AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_1934_), .C(_1905_), .D(_1913_), .Y(_2123_) );
	OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2122_), .B(_2123_), .C(_1930_), .Y(_2124_) );
	XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2124_), .B(_2118_), .Y(_2125_) );
	NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(divider_divuResult_18_bF_buf1), .Y(_2126_) );
	NAND3X1 NAND3X1_433 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_2126_), .C(_2117_), .Y(_2127_) );
	INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .Y(_2128_) );
	NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(divider_divuResult_18_bF_buf0), .Y(_2129_) );
	AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf5), .B(_2125_), .Y(_2131_) );
	OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(_2131_), .C(_4999__bF_buf5), .Y(_2132_) );
	XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(_2122_), .Y(_2133_) );
	INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .Y(_2134_) );
	NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(divider_divuResult_18_bF_buf4), .Y(_2135_) );
	OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf3), .B(_1983__bF_buf4), .C(_2120_), .Y(_2136_) );
	NAND3X1 NAND3X1_434 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_2135_), .C(_2136_), .Y(_2137_) );
	NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(divider_divuResult_18_bF_buf3), .Y(_2138_) );
	OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf2), .B(_1983__bF_buf3), .C(_1939_), .Y(_2139_) );
	NAND3X1 NAND3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf3), .B(_2138_), .C(_2139_), .Y(_2140_) );
	AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(_2140_), .C(_2127_), .D(_2132_), .Y(_2142_) );
	OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf1), .B(_1983__bF_buf2), .C(_1923_), .Y(_2143_) );
	NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .B(_1894_), .Y(_2144_) );
	AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .B(_1904_), .Y(_2145_) );
	OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_19_), .B(divider_divuResult_19_bF_buf5), .C(_1908_), .Y(_2146_) );
	NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .B(_2146_), .Y(_2147_) );
	INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .Y(_2148_) );
	NAND3X1 NAND3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_2148_), .C(_2147_), .Y(_2149_) );
	AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_1910_), .C(_2145_), .Y(_2150_) );
	OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_1966_), .Y(_2151_) );
	AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(_2144_), .Y(_2153_) );
	NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2144_), .B(_2151_), .Y(_2154_) );
	OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(_2154_), .C(divider_divuResult_18_bF_buf2), .Y(_2155_) );
	NAND3X1 NAND3X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_2155_), .C(_2143_), .Y(_2156_) );
	INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .Y(_2157_) );
	NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1913_), .B(_2157_), .Y(_2158_) );
	OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2158_), .C(divider_divuResult_18_bF_buf1), .Y(_2159_) );
	OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf0), .B(_1983__bF_buf1), .C(_1932_), .Y(_2160_) );
	NAND3X1 NAND3X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf7), .B(_2159_), .C(_2160_), .Y(_2161_) );
	AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2155_), .C(_1735__bF_buf7), .Y(_2162_) );
	OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2161_), .B(_2162_), .C(_2156_), .Y(_2164_) );
	AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .B(_2126_), .C(_4999__bF_buf4), .Y(_2165_) );
	NAND3X1 NAND3X1_439 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf3), .B(_2126_), .C(_2117_), .Y(_2166_) );
	NAND3X1 NAND3X1_440 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_2135_), .C(_2136_), .Y(_2167_) );
	OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2165_), .C(_2166_), .Y(_2168_) );
	AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2164_), .B(_2142_), .C(_2168_), .Y(_2169_) );
	NAND3X1 NAND3X1_441 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .B(_2155_), .C(_2143_), .Y(_2170_) );
	INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .Y(_2171_) );
	OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf4), .B(_1983__bF_buf0), .C(_2171_), .Y(_2172_) );
	OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .B(_2150_), .C(_2144_), .Y(_2173_) );
	OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(_2144_), .Y(_2175_) );
	NAND3X1 NAND3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_2173_), .B(_2175_), .C(divider_divuResult_18_bF_buf0), .Y(_2176_) );
	NAND3X1 NAND3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf6), .B(_2176_), .C(_2172_), .Y(_2177_) );
	NAND3X1 NAND3X1_444 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .B(_2159_), .C(_2160_), .Y(_2178_) );
	NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2158_), .Y(_2179_) );
	NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .B(divider_divuResult_18_bF_buf5), .Y(_2180_) );
	INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .Y(_2181_) );
	OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf3), .B(_1983__bF_buf4), .C(_2181_), .Y(_2182_) );
	NAND3X1 NAND3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_2180_), .C(_2182_), .Y(_2183_) );
	AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2178_), .B(_2183_), .C(_2170_), .D(_2177_), .Y(_2184_) );
	NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_2184_), .B(_2142_), .Y(_2186_) );
	NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_2147_), .Y(_2187_) );
	XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_2187_), .B(_2148_), .Y(_2188_) );
	INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .Y(_2189_) );
	NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2189_), .B(divider_divuResult_18_bF_buf4), .Y(_2190_) );
	OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf2), .B(_1983__bF_buf3), .C(_2146_), .Y(_2191_) );
	AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2191_), .B(_2190_), .C(_2547__bF_buf1), .Y(_2192_) );
	INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_18_), .Y(_2193_) );
	NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf5), .B(_2193_), .Y(_2194_) );
	NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf0), .B(divider_aOp_abs_18_), .Y(_2195_) );
	OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2194_), .B(_2195_), .C(divider_divuResult_18_bF_buf3), .Y(_2197_) );
	OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf1), .B(_1983__bF_buf2), .C(_2193_), .Y(_2198_) );
	NAND3X1 NAND3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_2197_), .C(_2198_), .Y(_2199_) );
	NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .B(divider_divuResult_18_bF_buf2), .Y(_2200_) );
	OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2146_), .B(divider_divuResult_18_bF_buf1), .C(_2200_), .Y(_2201_) );
	NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_2201_), .Y(_2202_) );
	OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2199_), .B(_2192_), .C(_2202_), .Y(_2203_) );
	NAND3X1 NAND3X1_447 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_2197_), .C(_2198_), .Y(_2204_) );
	NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .B(_2193_), .Y(_2205_) );
	OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_2205_), .C(divider_divuResult_18_bF_buf0), .Y(_2206_) );
	OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf0), .B(_1983__bF_buf1), .C(divider_aOp_abs_18_), .Y(_2208_) );
	NAND3X1 NAND3X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf2), .B(_2206_), .C(_2208_), .Y(_2209_) );
	NAND3X1 NAND3X1_449 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_2190_), .C(_2191_), .Y(_2210_) );
	INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(_2146_), .Y(_2211_) );
	OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_1699__bF_buf4), .B(_1983__bF_buf0), .C(_2211_), .Y(_2212_) );
	NAND3X1 NAND3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_2200_), .C(_2212_), .Y(_2213_) );
	AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2209_), .C(_2210_), .D(_2213_), .Y(_2214_) );
	NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_17_), .B(_1746__bF_buf4), .Y(_2215_) );
	INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .Y(_2216_) );
	INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_17_), .Y(_2217_) );
	NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_2217_), .Y(_2219_) );
	AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2216_), .B(divider_aOp_abs_16_), .C(_2219_), .Y(_2220_) );
	INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(_2220_), .Y(_2221_) );
	AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2221_), .C(_2203_), .Y(_2222_) );
	OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2222_), .C(_2169_), .Y(_2223_) );
	NAND3X1 NAND3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .B(_2116_), .C(_2223_), .Y(_2224_) );
	INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_16_), .Y(_2225_) );
	NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .B(_2219_), .Y(_2226_) );
	NAND3X1 NAND3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_2226_), .C(_2214_), .Y(_2227_) );
	NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2227_), .Y(_2228_) );
	NAND3X1 NAND3X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2033_), .C(_2228_), .Y(_2230_) );
	NAND3X1 NAND3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2106_), .B(_2230_), .C(_2224_), .Y(_2231_) );
	AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .B(_1946_), .C(_1948_), .Y(_2232_) );
	OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf1), .B(_2232_), .C(_1944__bF_buf4), .Y(_2233_) );
	NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_2164_), .Y(_2234_) );
	INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(_2168_), .Y(_2235_) );
	NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(_2234_), .Y(_2236_) );
	INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .Y(_2237_) );
	OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2211_), .B(divider_divuResult_18_bF_buf5), .C(_2190_), .Y(_2238_) );
	NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_2238_), .Y(_2239_) );
	INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(_2199_), .Y(_2241_) );
	NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_2238_), .Y(_2242_) );
	AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_2241_), .B(_2239_), .C(_2242_), .Y(_2243_) );
	AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2206_), .C(_1768__bF_buf1), .Y(_2244_) );
	AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .B(_2197_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .Y(_2245_) );
	AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2212_), .B(_2200_), .C(_2547__bF_buf6), .Y(_2246_) );
	AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2191_), .B(_2190_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .Y(_2247_) );
	OAI22X1 OAI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .B(_2245_), .C(_2246_), .D(_2247_), .Y(_2248_) );
	OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2248_), .B(_2220_), .C(_2243_), .Y(_2249_) );
	AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_2249_), .C(_2236_), .Y(_2250_) );
	NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2033_), .Y(_2252_) );
	OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .B(_2250_), .C(_2106_), .Y(_2253_) );
	INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(_2230_), .Y(_2254_) );
	OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_2254_), .B(_2253_), .C(_1946_), .Y(_2255_) );
	NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(_2255__bF_buf4), .Y(_2256_) );
	NAND3X1 NAND3X1_455 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .B(_2229__bF_buf4), .C(_2256_), .Y(_2257_) );
	AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_2257_), .B(_2233_), .Y(_2258_) );
	INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .Y(_2259_) );
	OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_2074_), .B(_2115_), .Y(_2260_) );
	NAND3X1 NAND3X1_456 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .B(_2206_), .C(_2208_), .Y(_2261_) );
	NAND3X1 NAND3X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2216_), .B(_2199_), .C(_2261_), .Y(_2263_) );
	OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(divider_divuResult_18_bF_buf4), .C(_2206_), .Y(_2264_) );
	AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2201_), .B(_2547__bF_buf5), .C(_1768__bF_buf0), .D(_2264_), .Y(_2265_) );
	AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .B(_2238_), .C(_2265_), .D(_2263_), .Y(_2266_) );
	NAND3X1 NAND3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_2184_), .C(_2266_), .Y(_2267_) );
	AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2169_), .C(_2260_), .Y(_2268_) );
	OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2268_), .C(_2033_), .Y(_2269_) );
	AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_2259_), .C(_1945_), .Y(divider_divuResult_17_) );
	NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1985_), .Y(_2270_) );
	INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .Y(_2271_) );
	OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2268_), .C(_2271_), .Y(_2273_) );
	AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_2013_), .C(_2270_), .Y(_2274_) );
	INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(_2270_), .Y(_2275_) );
	AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2209_), .C(_2215_), .Y(_2276_) );
	OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_2238_), .C(_2199_), .Y(_2277_) );
	OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_2277_), .B(_2276_), .C(_2239_), .Y(_2278_) );
	OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2278_), .C(_2169_), .Y(_2279_) );
	AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2116_), .C(_2105_), .Y(_2280_) );
	OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_2280_), .C(_2013_), .Y(_2281_) );
	NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_2281_), .Y(_2282_) );
	OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_2274_), .B(_2282_), .C(divider_divuResult_17_bF_buf3), .Y(_2284_) );
	OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_1951_), .B(divider_divuResult_18_bF_buf3), .C(_1982_), .Y(_2285_) );
	NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(_2255__bF_buf3), .Y(_2286_) );
	NAND3X1 NAND3X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf3), .B(_2286_), .C(_2284_), .Y(_2287_) );
	NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_2281_), .Y(_2288_) );
	NAND3X1 NAND3X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2270_), .B(_2013_), .C(_2273_), .Y(_2289_) );
	NAND3X1 NAND3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2289_), .B(_2288_), .C(divider_divuResult_17_bF_buf2), .Y(_2290_) );
	NAND3X1 NAND3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_1984_), .C(_2255__bF_buf2), .Y(_2291_) );
	NAND3X1 NAND3X1_463 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf1), .B(_2291_), .C(_2290_), .Y(_2292_) );
	NAND3X1 NAND3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2287_), .B(_2292_), .C(_2258_), .Y(_2293_) );
	OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_2003_), .B(divider_divuResult_18_bF_buf2), .C(_2023_), .Y(_2295_) );
	NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .B(_2255__bF_buf1), .Y(_2296_) );
	INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .Y(_2297_) );
	NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2006_), .Y(_2298_) );
	INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(_2298_), .Y(_2299_) );
	OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2268_), .C(_2030_), .Y(_2300_) );
	NAND3X1 NAND3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2297_), .B(_2299_), .C(_2300_), .Y(_2301_) );
	INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .Y(_2302_) );
	INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .Y(_2303_) );
	NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2279_), .Y(_2304_) );
	AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .B(_2303_), .C(_2302_), .Y(_2306_) );
	OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2306_), .C(_2298_), .Y(_2307_) );
	NAND3X1 NAND3X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2301_), .B(_2307_), .C(divider_divuResult_17_bF_buf1), .Y(_2308_) );
	NAND3X1 NAND3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf1), .B(_2296_), .C(_2308_), .Y(_2309_) );
	OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2306_), .C(_2299_), .Y(_2310_) );
	NAND3X1 NAND3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2297_), .B(_2298_), .C(_2300_), .Y(_2311_) );
	NAND3X1 NAND3X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2311_), .B(_2310_), .C(divider_divuResult_17_bF_buf0), .Y(_2312_) );
	INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .Y(_2313_) );
	NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(_2255__bF_buf0), .Y(_2314_) );
	NAND3X1 NAND3X1_470 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_2314_), .C(_2312_), .Y(_2315_) );
	NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2280_), .Y(_2317_) );
	NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .B(_2317_), .Y(_2318_) );
	NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .B(divider_divuResult_17_bF_buf3), .Y(_2319_) );
	NAND3X1 NAND3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(_2011_), .C(_2255__bF_buf4), .Y(_2320_) );
	NAND3X1 NAND3X1_472 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .B(_2320_), .C(_2319_), .Y(_2321_) );
	OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_2255__bF_buf3), .B(_2318_), .Y(_2322_) );
	NAND3X1 NAND3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(_2027_), .C(_2255__bF_buf2), .Y(_2323_) );
	NAND3X1 NAND3X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf0), .B(_2323_), .C(_2322_), .Y(_2324_) );
	NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2321_), .B(_2324_), .Y(_2325_) );
	NAND3X1 NAND3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_2309_), .B(_2315_), .C(_2325_), .Y(_2326_) );
	NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2326_), .Y(_2328_) );
	OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(divider_divuResult_18_bF_buf1), .C(_2050_), .Y(_2329_) );
	NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2329_), .B(_2255__bF_buf1), .Y(_2330_) );
	NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2051_), .B(_2058_), .Y(_2331_) );
	INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .Y(_2332_) );
	INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(_2103_), .Y(_2333_) );
	INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2334_) );
	AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2169_), .C(_2115_), .Y(_2335_) );
	OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2335_), .C(_2073_), .Y(_2336_) );
	NAND3X1 NAND3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .B(_2333_), .C(_2336_), .Y(_2337_) );
	INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(_2073_), .Y(_2339_) );
	INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2340_) );
	OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_2088_), .C(_2340_), .Y(_2341_) );
	INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .Y(_2342_) );
	AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .B(_2341_), .C(_2342_), .D(_2279_), .Y(_2343_) );
	OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2343_), .C(_2333_), .Y(_2344_) );
	NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .B(_2344_), .Y(_2345_) );
	NAND3X1 NAND3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2337_), .B(_2345_), .C(divider_divuResult_17_bF_buf2), .Y(_2346_) );
	NAND3X1 NAND3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf4), .B(_2330_), .C(_2346_), .Y(_2347_) );
	NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .B(_2344_), .Y(_2348_) );
	NAND3X1 NAND3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .B(_2333_), .C(_2336_), .Y(_2350_) );
	NAND3X1 NAND3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2350_), .B(_2348_), .C(divider_divuResult_17_bF_buf1), .Y(_2351_) );
	INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(_2329_), .Y(_2352_) );
	NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2352_), .B(_2255__bF_buf0), .Y(_2353_) );
	NAND3X1 NAND3X1_481 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .B(_2353_), .C(_2351_), .Y(_2354_) );
	AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_2347_), .B(_2354_), .Y(_2355_) );
	NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .B(_2343_), .Y(_2356_) );
	NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_2356_), .B(_2336_), .Y(_2357_) );
	NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2357_), .B(divider_divuResult_17_bF_buf0), .Y(_2358_) );
	NAND3X1 NAND3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2069_), .B(_2071_), .C(_2255__bF_buf4), .Y(_2359_) );
	NAND3X1 NAND3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf4), .B(_2359_), .C(_2358_), .Y(_2361_) );
	AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_2336_), .B(_2356_), .Y(_2362_) );
	NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2362_), .B(divider_divuResult_17_bF_buf3), .Y(_2363_) );
	NAND3X1 NAND3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2066_), .C(_2255__bF_buf3), .Y(_2364_) );
	NAND3X1 NAND3X1_485 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .B(_2364_), .C(_2363_), .Y(_2365_) );
	AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .B(_2365_), .Y(_2366_) );
	NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2366_), .B(_2355_), .Y(_2367_) );
	NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_2110_), .Y(_2368_) );
	INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(_2368_), .Y(_2369_) );
	NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2114_), .Y(_2370_) );
	AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2169_), .C(_2370_), .Y(_2372_) );
	OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .B(_2372_), .C(_2369_), .Y(_2373_) );
	OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2114_), .C(_2279_), .Y(_2374_) );
	NAND3X1 NAND3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2368_), .C(_2374_), .Y(_2375_) );
	AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .B(_2375_), .Y(_2376_) );
	NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2255__bF_buf2), .Y(_2377_) );
	OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_2255__bF_buf1), .B(_2376_), .C(_2377_), .Y(_2378_) );
	NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .B(_2378_), .Y(_2379_) );
	NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .B(_2378_), .Y(_2380_) );
	OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(divider_divuResult_18_bF_buf0), .C(_2099_), .Y(_2381_) );
	NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2381_), .B(_2255__bF_buf0), .Y(_2383_) );
	XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2370_), .Y(_2384_) );
	NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2384_), .B(divider_divuResult_17_bF_buf2), .Y(_2385_) );
	AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2385_), .B(_2383_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .Y(_2386_) );
	OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_2386_), .B(_2380_), .C(_2379_), .Y(_2387_) );
	INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(_2347_), .Y(_2388_) );
	INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .Y(_2389_) );
	AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_2354_), .C(_2388_), .Y(_2390_) );
	OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .B(_2367_), .C(_2390_), .Y(_2391_) );
	OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(divider_divuResult_17_bF_buf1), .C(_2308_), .Y(_2392_) );
	INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .Y(_2394_) );
	OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_2255__bF_buf4), .B(_2318_), .C(_2323_), .Y(_2395_) );
	NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf4), .B(_2395_), .Y(_2396_) );
	OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .B(_2392_), .C(_2396_), .Y(_2397_) );
	OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf0), .B(_2394_), .C(_2397_), .Y(_2398_) );
	NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2233_), .B(_2257_), .Y(_2399_) );
	OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .B(_2287_), .C(_2233_), .Y(_2400_) );
	INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .Y(_2401_) );
	OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2398_), .C(_2401_), .Y(_2402_) );
	AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_2328_), .C(_2402_), .Y(_2403_) );
	OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(_2131_), .C(_2255__bF_buf3), .Y(_2405_) );
	NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(_2132_), .Y(_2406_) );
	INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .Y(_2407_) );
	INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(_2164_), .Y(_2408_) );
	NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2184_), .B(_2266_), .Y(_2409_) );
	AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(_2140_), .C(_2408_), .D(_2409_), .Y(_2410_) );
	OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_2407_), .B(_2410_), .C(_2406_), .Y(_2411_) );
	INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(_2406_), .Y(_2412_) );
	NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(_2140_), .Y(_2413_) );
	NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .B(_2409_), .Y(_2414_) );
	NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(_2414_), .Y(_2416_) );
	NAND3X1 NAND3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2412_), .B(_2167_), .C(_2416_), .Y(_2417_) );
	NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2411_), .B(_2417_), .Y(_2418_) );
	NAND3X1 NAND3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2231_), .C(_2418_), .Y(_2419_) );
	NAND3X1 NAND3X1_489 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .B(_2405_), .C(_2419_), .Y(_2420_) );
	OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(divider_divuResult_18_bF_buf5), .C(_2126_), .Y(_2421_) );
	INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .Y(_2422_) );
	AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .B(_1946_), .C(_2422_), .Y(_2423_) );
	AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2411_), .B(_2417_), .C(_2255__bF_buf2), .Y(_2424_) );
	OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2424_), .C(_4714__bF_buf5), .Y(_2425_) );
	NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(_2414_), .Y(_2427_) );
	OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(_2410_), .Y(_2428_) );
	NAND3X1 NAND3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2231_), .C(_2428_), .Y(_2429_) );
	OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_1939_), .B(divider_divuResult_18_bF_buf4), .C(_2135_), .Y(_2430_) );
	NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .B(_2255__bF_buf1), .Y(_2431_) );
	NAND3X1 NAND3X1_491 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .B(_2429_), .C(_2431_), .Y(_2432_) );
	NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .B(_2427_), .Y(_2433_) );
	NAND3X1 NAND3X1_492 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2231_), .C(_2433_), .Y(_2434_) );
	INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .Y(_2435_) );
	NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2435_), .B(_2255__bF_buf0), .Y(_2436_) );
	NAND3X1 NAND3X1_493 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf2), .B(_2434_), .C(_2436_), .Y(_2438_) );
	AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .B(_2438_), .C(_2420_), .D(_2425_), .Y(_2439_) );
	OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(divider_divuResult_18_bF_buf3), .C(_2155_), .Y(_2440_) );
	NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2440_), .B(_2255__bF_buf4), .Y(_2441_) );
	NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2170_), .B(_2177_), .Y(_2442_) );
	NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2178_), .B(_2183_), .Y(_2443_) );
	INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .Y(_2444_) );
	OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(_2278_), .C(_2161_), .Y(_2445_) );
	XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2445_), .B(_2442_), .Y(_2446_) );
	NAND3X1 NAND3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2446_), .C(_2231_), .Y(_2447_) );
	NAND3X1 NAND3X1_495 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .B(_2447_), .C(_2441_), .Y(_2449_) );
	INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(_2440_), .Y(_2450_) );
	NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(_2255__bF_buf3), .Y(_2451_) );
	INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .Y(_2452_) );
	NAND3X1 NAND3X1_496 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2231_), .C(_2452_), .Y(_2453_) );
	NAND3X1 NAND3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf1), .B(_2453_), .C(_2451_), .Y(_2454_) );
	XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2266_), .B(_2444_), .Y(_2455_) );
	INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .Y(_2456_) );
	NAND3X1 NAND3X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2456_), .C(_2231_), .Y(_2457_) );
	OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_2181_), .B(divider_divuResult_18_bF_buf2), .C(_2159_), .Y(_2458_) );
	NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2458_), .B(_2255__bF_buf2), .Y(_2460_) );
	NAND3X1 NAND3X1_499 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .B(_2457_), .C(_2460_), .Y(_2461_) );
	NAND3X1 NAND3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2455_), .C(_2231_), .Y(_2462_) );
	INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(_2458_), .Y(_2463_) );
	NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_2255__bF_buf1), .Y(_2464_) );
	NAND3X1 NAND3X1_501 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf5), .B(_2462_), .C(_2464_), .Y(_2465_) );
	AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2454_), .C(_2461_), .D(_2465_), .Y(_2466_) );
	NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_2439_), .Y(_2467_) );
	NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_2210_), .B(_2213_), .Y(_2468_) );
	INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(_2261_), .Y(_2469_) );
	OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .B(_2469_), .C(_2199_), .Y(_2471_) );
	XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .B(_2468_), .Y(_2472_) );
	NAND3X1 NAND3X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2472_), .C(_2231_), .Y(_2473_) );
	NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2238_), .B(_2255__bF_buf0), .Y(_2474_) );
	NAND3X1 NAND3X1_503 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_2473_), .C(_2474_), .Y(_2475_) );
	INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .Y(_2476_) );
	AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .B(_1946_), .C(_2201_), .Y(_2477_) );
	OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2476_), .C(_2470__bF_buf5), .Y(_2478_) );
	OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_2241_), .B(_2469_), .C(_2215_), .Y(_2479_) );
	NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2263_), .B(_2479_), .Y(_2480_) );
	NAND3X1 NAND3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2480_), .C(_2231_), .Y(_2482_) );
	OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_18_), .B(divider_divuResult_18_bF_buf1), .C(_2197_), .Y(_2483_) );
	NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .B(_2255__bF_buf4), .Y(_2484_) );
	NAND3X1 NAND3X1_505 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_2482_), .C(_2484_), .Y(_2485_) );
	NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .B(_2255__bF_buf3), .Y(_2486_) );
	INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(_2480_), .Y(_2487_) );
	NAND3X1 NAND3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2487_), .C(_2231_), .Y(_2488_) );
	NAND3X1 NAND3X1_507 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_2488_), .C(_2486_), .Y(_2489_) );
	AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_2485_), .B(_2489_), .C(_2475_), .D(_2478_), .Y(_2490_) );
	NAND3X1 NAND3X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2226_), .C(_2231_), .Y(_2491_) );
	NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2217_), .B(_2255__bF_buf2), .Y(_2493_) );
	AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2493_), .B(_2491_), .C(_1768__bF_buf7), .Y(_2494_) );
	NAND3X1 NAND3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf6), .B(_2491_), .C(_2493_), .Y(_2495_) );
	NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(_2225_), .Y(_2496_) );
	INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .Y(_2497_) );
	AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .B(_2497_), .C(_2494_), .Y(_2498_) );
	NAND3X1 NAND3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf4), .B(_2473_), .C(_2474_), .Y(_2499_) );
	AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2473_), .C(_2470__bF_buf3), .Y(_2500_) );
	NAND3X1 NAND3X1_511 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_2482_), .C(_2484_), .Y(_2501_) );
	OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .B(_2500_), .C(_2499_), .Y(_2502_) );
	AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2490_), .B(_2498_), .C(_2502_), .Y(_2504_) );
	NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(_2504_), .Y(_2505_) );
	AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2441_), .B(_2447_), .C(_4100__bF_buf0), .Y(_2506_) );
	NAND3X1 NAND3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf7), .B(_2447_), .C(_2441_), .Y(_2507_) );
	NAND3X1 NAND3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf4), .B(_2457_), .C(_2460_), .Y(_2508_) );
	AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .B(_2508_), .C(_2506_), .Y(_2509_) );
	NAND3X1 NAND3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf4), .B(_2405_), .C(_2419_), .Y(_2510_) );
	AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2419_), .B(_2405_), .C(_4714__bF_buf3), .Y(_2511_) );
	NAND3X1 NAND3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_2429_), .C(_2431_), .Y(_2512_) );
	OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_2512_), .B(_2511_), .C(_2510_), .Y(_2513_) );
	AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2439_), .B(_2509_), .C(_2513_), .Y(_2515_) );
	NAND3X1 NAND3X1_516 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .B(_2491_), .C(_2493_), .Y(_2516_) );
	INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(_2226_), .Y(_2517_) );
	NAND3X1 NAND3X1_517 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_2517_), .C(_2231_), .Y(_2518_) );
	NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_17_), .B(_2255__bF_buf1), .Y(_2519_) );
	NAND3X1 NAND3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_2518_), .C(_2519_), .Y(_2520_) );
	NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(divider_aOp_abs_16_), .Y(_2521_) );
	NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf3), .B(_2225_), .Y(_2522_) );
	NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .B(_2522_), .Y(_2523_) );
	INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .Y(_2524_) );
	AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2516_), .B(_2520_), .C(_2524_), .Y(_2526_) );
	NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .B(_2490_), .Y(_2527_) );
	OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(_2527_), .C(_2515_), .Y(_2528_) );
	NAND3X1 NAND3X1_519 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf0), .B(_2286_), .C(_2284_), .Y(_2529_) );
	NAND3X1 NAND3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf2), .B(_2291_), .C(_2290_), .Y(_2530_) );
	AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .B(_2530_), .C(_2399_), .Y(_2531_) );
	AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_2309_), .B(_2315_), .Y(_2532_) );
	NAND3X1 NAND3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .B(_2325_), .C(_2531_), .Y(_2533_) );
	NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2375_), .B(_2373_), .Y(_2534_) );
	NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2534_), .B(divider_divuResult_17_bF_buf0), .Y(_2535_) );
	NAND3X1 NAND3X1_522 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_2377_), .C(_2535_), .Y(_2537_) );
	NAND3X1 NAND3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2087_), .C(_2255__bF_buf0), .Y(_2538_) );
	NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_2376_), .B(divider_divuResult_17_bF_buf3), .Y(_2539_) );
	NAND3X1 NAND3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf0), .B(_2538_), .C(_2539_), .Y(_2540_) );
	OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_2255__bF_buf4), .B(_2384_), .Y(_2541_) );
	INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(_2381_), .Y(_2542_) );
	NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2542_), .B(_2255__bF_buf3), .Y(_2543_) );
	NAND3X1 NAND3X1_525 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .B(_2543_), .C(_2541_), .Y(_2544_) );
	NAND3X1 NAND3X1_526 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf0), .B(_2383_), .C(_2385_), .Y(_2545_) );
	AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .B(_2540_), .C(_2545_), .D(_2544_), .Y(_2546_) );
	NAND3X1 NAND3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2366_), .B(_2546_), .C(_2355_), .Y(_2548_) );
	NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2548_), .B(_2533_), .Y(_2549_) );
	OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .B(_2528_), .C(_2549_), .Y(_2550_) );
	AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2403_), .C(_3204__bF_buf3), .Y(divider_divuResult_16_) );
	OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_2256_), .B(divider_divuResult_16_bF_buf5), .C(_2229__bF_buf3), .Y(_2551_) );
	XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(divider_absoluteValue_B_flipSign_result_16_bF_buf3), .Y(_2552_) );
	INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(_2326_), .Y(_2553_) );
	AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_2439_), .B(_2466_), .Y(_2554_) );
	NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_2477_), .C(_2476_), .Y(_2555_) );
	AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2473_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .Y(_2556_) );
	AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(_2488_), .C(_2547__bF_buf2), .Y(_2558_) );
	AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2484_), .B(_2482_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .Y(_2559_) );
	OAI22X1 OAI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_2558_), .B(_2559_), .C(_2556_), .D(_2555_), .Y(_2560_) );
	OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_17_), .B(divider_divuResult_17_bF_buf2), .C(_2491_), .Y(_2561_) );
	NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_2561_), .Y(_2562_) );
	AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2519_), .B(_2518_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .Y(_2563_) );
	OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .B(_2563_), .C(_2562_), .Y(_2564_) );
	INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .Y(_2565_) );
	OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2476_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .Y(_2566_) );
	AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(_2488_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .Y(_2567_) );
	AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2567_), .C(_2565_), .Y(_2569_) );
	OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_2564_), .B(_2560_), .C(_2569_), .Y(_2570_) );
	NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(_2570_), .Y(_2571_) );
	NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf2), .B(_2423_), .C(_2424_), .Y(_2572_) );
	AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2419_), .B(_2405_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .Y(_2573_) );
	NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .B(_2438_), .Y(_2574_) );
	OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .B(_2572_), .C(_2574_), .Y(_2575_) );
	OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(divider_divuResult_17_bF_buf1), .C(_2447_), .Y(_2576_) );
	NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .B(_2576_), .Y(_2577_) );
	AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2453_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .Y(_2578_) );
	AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2462_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .Y(_2580_) );
	OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2580_), .C(_2577_), .Y(_2581_) );
	INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(_2510_), .Y(_2582_) );
	OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2424_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .Y(_2583_) );
	INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(_2512_), .Y(_2584_) );
	AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_2583_), .C(_2582_), .Y(_2585_) );
	OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .B(_2575_), .C(_2585_), .Y(_2586_) );
	AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_2490_), .B(_2526_), .Y(_2587_) );
	AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(_2587_), .C(_2586_), .Y(_2588_) );
	AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2571_), .C(_2548_), .Y(_2589_) );
	OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_2589_), .C(_2553_), .Y(_2591_) );
	AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .B(_2530_), .C(_2398_), .D(_2591_), .Y(_2592_) );
	NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2530_), .B(_2529_), .Y(_2593_) );
	NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_2309_), .B(_2315_), .Y(_2594_) );
	OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_2396_), .B(_2594_), .C(_2309_), .Y(_2595_) );
	NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2347_), .B(_2354_), .Y(_2596_) );
	NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .B(_2365_), .Y(_2597_) );
	NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_2596_), .Y(_2598_) );
	OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_2255__bF_buf2), .B(_2534_), .C(_2538_), .Y(_2599_) );
	NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf6), .B(_2599_), .Y(_2600_) );
	NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf5), .B(_2599_), .Y(_2602_) );
	OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_2542_), .B(divider_divuResult_17_bF_buf0), .C(_2385_), .Y(_2603_) );
	NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf5), .B(_2603_), .Y(_2604_) );
	AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2604_), .B(_2602_), .C(_2600_), .Y(_2605_) );
	OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .B(_2596_), .C(_2347_), .Y(_2606_) );
	AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2598_), .B(_2605_), .C(_2606_), .Y(_2607_) );
	INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(_2548_), .Y(_2608_) );
	OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .B(_2528_), .C(_2608_), .Y(_2609_) );
	AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2609_), .B(_2607_), .C(_2326_), .Y(_2610_) );
	NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_2593_), .B(_2595_), .C(_2610_), .Y(_2611_) );
	OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_2611_), .B(_2592_), .C(divider_divuResult_16_bF_buf4), .Y(_2613_) );
	OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(divider_divuResult_17_bF_buf3), .C(_2290_), .Y(_2614_) );
	INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(_2614_), .Y(_2615_) );
	AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(_2531_), .C(_2400_), .Y(_2616_) );
	OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .B(_2607_), .C(_2616_), .Y(_2617_) );
	NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_2554_), .Y(_2618_) );
	NAND3X1 NAND3X1_528 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .B(_2618_), .C(_2571_), .Y(_2619_) );
	AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2549_), .C(_2617_), .Y(_2620_) );
	OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf2), .B(_2620__bF_buf4), .C(_2615_), .Y(_2621_) );
	NAND3X1 NAND3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf3), .B(_2621_), .C(_2613_), .Y(_2622_) );
	OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf1), .B(_2620__bF_buf3), .C(_2614_), .Y(_2624_) );
	OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(_2610_), .C(_2593_), .Y(_2625_) );
	INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(_2593_), .Y(_2626_) );
	NAND3X1 NAND3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .B(_2398_), .C(_2591_), .Y(_2627_) );
	NAND3X1 NAND3X1_531 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf3), .B(_2625_), .C(_2627_), .Y(_2628_) );
	NAND3X1 NAND3X1_532 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .B(_2624_), .C(_2628_), .Y(_2629_) );
	NAND3X1 NAND3X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .B(_2629_), .C(_2622_), .Y(_2630_) );
	OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf0), .B(_2620__bF_buf2), .C(_2392_), .Y(_2631_) );
	OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_2589_), .C(_2325_), .Y(_2632_) );
	NAND3X1 NAND3X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .B(_2396_), .C(_2632_), .Y(_2633_) );
	INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(_2396_), .Y(_2635_) );
	INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(_2325_), .Y(_2636_) );
	AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2609_), .B(_2607_), .C(_2636_), .Y(_2637_) );
	OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2637_), .C(_2594_), .Y(_2638_) );
	NAND3X1 NAND3X1_535 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf2), .B(_2638_), .C(_2633_), .Y(_2639_) );
	NAND3X1 NAND3X1_536 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf1), .B(_2631_), .C(_2639_), .Y(_2640_) );
	OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf4), .B(_2620__bF_buf1), .C(_2394_), .Y(_2641_) );
	OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2637_), .C(_2532_), .Y(_2642_) );
	NAND3X1 NAND3X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2594_), .B(_2396_), .C(_2632_), .Y(_2643_) );
	NAND3X1 NAND3X1_538 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf1), .B(_2642_), .C(_2643_), .Y(_2644_) );
	NAND3X1 NAND3X1_539 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .B(_2641_), .C(_2644_), .Y(_2646_) );
	NAND3X1 NAND3X1_540 ( .gnd(gnd), .vdd(vdd), .A(_2636_), .B(_2607_), .C(_2609_), .Y(_2647_) );
	INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .Y(_2648_) );
	OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_2637_), .B(_2648_), .C(divider_divuResult_16_bF_buf0), .Y(_2649_) );
	INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(_2395_), .Y(_2650_) );
	OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf3), .B(_2620__bF_buf0), .C(_2650_), .Y(_2651_) );
	NAND3X1 NAND3X1_541 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .B(_2651_), .C(_2649_), .Y(_2652_) );
	OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf2), .B(_2620__bF_buf4), .C(_2395_), .Y(_2653_) );
	NAND3X1 NAND3X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .B(divider_divuResult_16_bF_buf5), .C(_2632_), .Y(_2654_) );
	NAND3X1 NAND3X1_543 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf4), .B(_2653_), .C(_2654_), .Y(_2655_) );
	NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2655_), .B(_2652_), .Y(_2657_) );
	NAND3X1 NAND3X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2646_), .C(_2657_), .Y(_2658_) );
	NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2630_), .Y(_2659_) );
	OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .B(_2528_), .C(_2546_), .Y(_2660_) );
	AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2660_), .B(_2387_), .C(_2597_), .Y(_2661_) );
	OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_2661_), .C(_2355_), .Y(_2662_) );
	AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .B(_2538_), .C(_8971__bF_buf4), .Y(_2663_) );
	AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .B(_2377_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .Y(_2664_) );
	AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2385_), .B(_2383_), .C(_7204__bF_buf4), .Y(_2665_) );
	AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .B(_2543_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .Y(_2666_) );
	OAI22X1 OAI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_2663_), .B(_2664_), .C(_2665_), .D(_2666_), .Y(_2668_) );
	AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2571_), .C(_2668_), .Y(_2669_) );
	OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .B(_2669_), .C(_2366_), .Y(_2670_) );
	NAND3X1 NAND3X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2596_), .B(_2361_), .C(_2670_), .Y(_2671_) );
	NAND3X1 NAND3X1_546 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf4), .B(_2662_), .C(_2671_), .Y(_2672_) );
	OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_2352_), .B(divider_divuResult_17_bF_buf2), .C(_2346_), .Y(_2673_) );
	INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .Y(_2674_) );
	OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf1), .B(_2620__bF_buf3), .C(_2674_), .Y(_2675_) );
	NAND3X1 NAND3X1_547 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .B(_2675_), .C(_2672_), .Y(_2676_) );
	AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2672_), .B(_2675_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .Y(_2677_) );
	OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_2255__bF_buf1), .B(_2362_), .C(_2359_), .Y(_2679_) );
	INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(_2679_), .Y(_2680_) );
	NAND3X1 NAND3X1_548 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_2387_), .C(_2660_), .Y(_2681_) );
	INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(_2681_), .Y(_2682_) );
	OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_2661_), .B(_2682_), .C(divider_divuResult_16_bF_buf3), .Y(_2683_) );
	OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_2680_), .B(divider_divuResult_16_bF_buf2), .C(_2683_), .Y(_2684_) );
	NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .B(_2684_), .Y(_2685_) );
	OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_2677_), .B(_2685_), .C(_2676_), .Y(_2686_) );
	OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf0), .B(_2620__bF_buf2), .C(_2673_), .Y(_2687_) );
	NAND3X1 NAND3X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2355_), .B(_2361_), .C(_2670_), .Y(_2688_) );
	OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_2661_), .C(_2596_), .Y(_2690_) );
	NAND3X1 NAND3X1_550 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf1), .B(_2690_), .C(_2688_), .Y(_2691_) );
	NAND3X1 NAND3X1_551 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf3), .B(_2687_), .C(_2691_), .Y(_2692_) );
	OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf4), .B(_2620__bF_buf1), .C(_2679_), .Y(_2693_) );
	NAND3X1 NAND3X1_552 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .B(_2693_), .C(_2683_), .Y(_2694_) );
	OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf3), .B(_2620__bF_buf0), .C(_2680_), .Y(_2695_) );
	NAND3X1 NAND3X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2681_), .B(divider_divuResult_16_bF_buf0), .C(_2670_), .Y(_2696_) );
	NAND3X1 NAND3X1_554 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf3), .B(_2695_), .C(_2696_), .Y(_2697_) );
	NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .B(_2694_), .Y(_2698_) );
	NAND3X1 NAND3X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2692_), .C(_2698_), .Y(_2699_) );
	NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2544_), .Y(_2701_) );
	AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2701_), .C(_2386_), .Y(_2702_) );
	OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_2663_), .B(_2664_), .C(_2702_), .Y(_2703_) );
	INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(_2603_), .Y(_2704_) );
	OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_2505_), .B(_2528_), .C(_2701_), .Y(_2705_) );
	OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .B(_2704_), .C(_2705_), .Y(_2706_) );
	OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_2600_), .B(_2380_), .C(_2706_), .Y(_2707_) );
	NAND3X1 NAND3X1_556 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf5), .B(_2707_), .C(_2703_), .Y(_2708_) );
	OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_2599_), .B(divider_divuResult_16_bF_buf4), .C(_2708_), .Y(_2709_) );
	NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .B(_2709_), .Y(_2710_) );
	OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf2), .B(_2620__bF_buf4), .C(_2599_), .Y(_2712_) );
	OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_2663_), .B(_2664_), .C(_2706_), .Y(_2713_) );
	OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_2600_), .B(_2380_), .C(_2702_), .Y(_2714_) );
	NAND3X1 NAND3X1_557 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf3), .B(_2713_), .C(_2714_), .Y(_2715_) );
	AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_2712_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .Y(_2716_) );
	OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf1), .B(_2620__bF_buf3), .C(_2603_), .Y(_2717_) );
	XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .B(_2701_), .Y(_2718_) );
	NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf2), .B(_2718_), .Y(_2719_) );
	AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2719_), .B(_2717_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .Y(_2720_) );
	OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_2720_), .B(_2716_), .C(_2710_), .Y(_2721_) );
	OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_2721_), .B(_2699_), .C(_2686_), .Y(_2723_) );
	AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(_2641_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .Y(_2724_) );
	AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_2654_), .B(_2653_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .Y(_2725_) );
	AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2646_), .B(_2725_), .C(_2724_), .Y(_2726_) );
	INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .Y(_2727_) );
	NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf2), .B(_2727_), .Y(_2728_) );
	AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2628_), .B(_2624_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .Y(_2729_) );
	AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2729_), .B(_2552_), .C(_2728_), .Y(_2730_) );
	OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_2726_), .B(_2630_), .C(_2730_), .Y(_2731_) );
	AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .B(_2659_), .C(_2731_), .Y(_2732_) );
	AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_2712_), .C(_10678__bF_buf3), .Y(_2734_) );
	OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf0), .B(_2620__bF_buf2), .C(_2378_), .Y(_2735_) );
	AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2708_), .B(_2735_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .Y(_2736_) );
	AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2719_), .B(_2717_), .C(_8971__bF_buf3), .Y(_2737_) );
	OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_2704_), .B(divider_divuResult_16_bF_buf1), .C(_2719_), .Y(_2738_) );
	NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .B(_2738_), .Y(_2739_) );
	OAI22X1 OAI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_2736_), .C(_2737_), .D(_2739_), .Y(_2740_) );
	NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .B(_2699_), .Y(_2741_) );
	AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .B(_2741_), .Y(_2742_) );
	AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2405_), .B(_2419_), .C(divider_divuResult_16_bF_buf0), .Y(_2743_) );
	INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf4), .Y(_2745_) );
	NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2608_), .B(_2328_), .Y(_2746_) );
	AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2571_), .C(_2746_), .Y(_2747_) );
	OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_2617_), .B(_2747_), .C(_2745_), .Y(_2748_) );
	NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2425_), .Y(_2749_) );
	INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2750_) );
	OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_2570_), .C(_2466_), .Y(_2751_) );
	AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2751_), .B(_2581_), .C(_2750_), .Y(_2752_) );
	OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_2752_), .C(_2749_), .Y(_2753_) );
	INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(_2749_), .Y(_2754_) );
	INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .Y(_2755_) );
	AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .B(_2527_), .C(_2755_), .Y(_2756_) );
	OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .B(_2756_), .C(_2574_), .Y(_2757_) );
	NAND3X1 NAND3X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2512_), .C(_2757_), .Y(_2758_) );
	AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_2758_), .C(_2748_), .Y(_2759_) );
	OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_2743_), .B(_2759_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .Y(_2760_) );
	OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_2422_), .B(divider_divuResult_17_bF_buf1), .C(_2419_), .Y(_2761_) );
	OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf3), .B(_2620__bF_buf1), .C(_2761_), .Y(_2762_) );
	NAND3X1 NAND3X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2749_), .B(_2512_), .C(_2757_), .Y(_2763_) );
	OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_2752_), .C(_2754_), .Y(_2764_) );
	NAND3X1 NAND3X1_560 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf5), .B(_2763_), .C(_2764_), .Y(_2766_) );
	NAND3X1 NAND3X1_561 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_2762_), .C(_2766_), .Y(_2767_) );
	OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .B(divider_divuResult_17_bF_buf0), .C(_2434_), .Y(_2768_) );
	NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2403_), .B(_2550_), .Y(_2769_) );
	NAND3X1 NAND3X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .B(_2581_), .C(_2751_), .Y(_2770_) );
	NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2770_), .B(_2757_), .Y(_2771_) );
	NAND3X1 NAND3X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2745_), .B(_2769_), .C(_2771_), .Y(_2772_) );
	OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(divider_divuResult_16_bF_buf4), .C(_2772_), .Y(_2773_) );
	OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .B(_2773_), .C(_2767_), .Y(_2774_) );
	NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_2774_), .Y(_2775_) );
	INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .Y(_2777_) );
	OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf2), .B(_2620__bF_buf0), .C(_2777_), .Y(_2778_) );
	NAND3X1 NAND3X1_564 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_2772_), .C(_2778_), .Y(_2779_) );
	AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_2757_), .B(_2770_), .Y(_2780_) );
	NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(divider_divuResult_16_bF_buf3), .Y(_2781_) );
	OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf1), .B(_2620__bF_buf4), .C(_2768_), .Y(_2782_) );
	NAND3X1 NAND3X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf1), .B(_2782_), .C(_2781_), .Y(_2783_) );
	NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_2779_), .B(_2783_), .Y(_2784_) );
	NAND3X1 NAND3X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_2767_), .C(_2784_), .Y(_2785_) );
	NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2454_), .Y(_2786_) );
	NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2465_), .Y(_2788_) );
	INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .Y(_2789_) );
	AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .B(_2527_), .C(_2789_), .Y(_2790_) );
	INVX1 INVX1_596 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .Y(_2791_) );
	NAND3X1 NAND3X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_2508_), .C(_2791_), .Y(_2792_) );
	INVX1 INVX1_597 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .Y(_2793_) );
	OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(_2790_), .C(_2793_), .Y(_2794_) );
	NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2794_), .B(_2792_), .Y(_2795_) );
	OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf0), .B(_2620__bF_buf3), .C(_2576_), .Y(_2796_) );
	OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2795_), .C(_2796_), .Y(_2797_) );
	NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_2797_), .Y(_2799_) );
	INVX1 INVX1_598 ( .gnd(gnd), .vdd(vdd), .A(_2576_), .Y(_2800_) );
	OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf4), .B(_2620__bF_buf2), .C(_2800_), .Y(_2801_) );
	NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf2), .B(_2795_), .Y(_2802_) );
	AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_2802_), .B(_2801_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .Y(_2803_) );
	OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(divider_divuResult_17_bF_buf3), .C(_2457_), .Y(_2804_) );
	INVX1 INVX1_599 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .Y(_2805_) );
	OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf3), .B(_2620__bF_buf1), .C(_2805_), .Y(_2806_) );
	INVX1 INVX1_600 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .Y(_2807_) );
	OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_2560_), .B(_2807_), .C(_2504_), .Y(_2808_) );
	NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_2808_), .Y(_2810_) );
	NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_2810_), .Y(_2811_) );
	NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_2811_), .B(divider_divuResult_16_bF_buf1), .Y(_2812_) );
	AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2812_), .B(_2806_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .Y(_2813_) );
	OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_2803_), .B(_2813_), .C(_2799_), .Y(_2814_) );
	OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .B(_2785_), .C(_2775_), .Y(_2815_) );
	INVX1 INVX1_601 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .Y(_2816_) );
	AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_2760_), .B(_2767_), .Y(_2817_) );
	NAND3X1 NAND3X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2792_), .B(_2794_), .C(divider_divuResult_16_bF_buf0), .Y(_2818_) );
	NAND3X1 NAND3X1_569 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .B(_2796_), .C(_2818_), .Y(_2819_) );
	NAND3X1 NAND3X1_570 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf0), .B(_2801_), .C(_2802_), .Y(_2821_) );
	OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_2810_), .C(divider_divuResult_16_bF_buf5), .Y(_2822_) );
	OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf2), .B(_2620__bF_buf0), .C(_2804_), .Y(_2823_) );
	NAND3X1 NAND3X1_571 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .B(_2823_), .C(_2822_), .Y(_2824_) );
	NAND3X1 NAND3X1_572 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf6), .B(_2806_), .C(_2812_), .Y(_2825_) );
	AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(_2825_), .C(_2819_), .D(_2821_), .Y(_2826_) );
	NAND3X1 NAND3X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2784_), .B(_2826_), .C(_2817_), .Y(_2827_) );
	NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2476_), .Y(_2828_) );
	OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf1), .B(_2620__bF_buf4), .C(_2828_), .Y(_2829_) );
	NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2478_), .Y(_2830_) );
	NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_2485_), .B(_2489_), .Y(_2832_) );
	OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .B(_2498_), .C(_2832_), .Y(_2833_) );
	INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(_2833_), .Y(_2834_) );
	OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_2567_), .B(_2834_), .C(_2830_), .Y(_2835_) );
	NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2567_), .B(_2834_), .Y(_2836_) );
	OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_2565_), .B(_2500_), .C(_2836_), .Y(_2837_) );
	NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_2835_), .B(_2837_), .Y(_2838_) );
	OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2838_), .C(_2829_), .Y(_2839_) );
	NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_2839_), .Y(_2840_) );
	INVX1 INVX1_602 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .Y(_2841_) );
	OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf0), .B(_2620__bF_buf3), .C(_2841_), .Y(_2843_) );
	NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_2838_), .B(divider_divuResult_16_bF_buf4), .Y(_2844_) );
	AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .B(_2843_), .C(_1735__bF_buf2), .Y(_2845_) );
	NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_2564_), .B(_2807_), .Y(_2846_) );
	NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2832_), .B(_2846_), .Y(_2847_) );
	OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2847_), .C(divider_divuResult_16_bF_buf3), .Y(_2848_) );
	OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .B(divider_divuResult_17_bF_buf2), .C(_2488_), .Y(_2849_) );
	INVX1 INVX1_603 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .Y(_2850_) );
	OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf4), .B(_2620__bF_buf2), .C(_2850_), .Y(_2851_) );
	NAND3X1 NAND3X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_2851_), .C(_2848_), .Y(_2852_) );
	OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_2845_), .B(_2852_), .C(_2840_), .Y(_2854_) );
	NAND3X1 NAND3X1_575 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .B(_2843_), .C(_2844_), .Y(_2855_) );
	AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_2837_), .B(_2835_), .Y(_2856_) );
	NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf2), .B(_2856_), .Y(_2857_) );
	NAND3X1 NAND3X1_576 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_2829_), .C(_2857_), .Y(_2858_) );
	NAND3X1 NAND3X1_577 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_2851_), .C(_2848_), .Y(_2859_) );
	NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2847_), .Y(_2860_) );
	NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_2860_), .B(divider_divuResult_16_bF_buf1), .Y(_2861_) );
	OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf3), .B(_2620__bF_buf1), .C(_2849_), .Y(_2862_) );
	NAND3X1 NAND3X1_578 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_2862_), .C(_2861_), .Y(_2863_) );
	AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_2858_), .C(_2859_), .D(_2863_), .Y(_2865_) );
	NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_2516_), .B(_2520_), .Y(_2866_) );
	NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_16_), .B(_1746__bF_buf2), .Y(_2867_) );
	XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_2866_), .B(_2867_), .Y(_2868_) );
	NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .B(divider_divuResult_16_bF_buf0), .Y(_2869_) );
	OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf2), .B(_2620__bF_buf0), .C(_2561_), .Y(_2870_) );
	NAND3X1 NAND3X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_2870_), .C(_2869_), .Y(_2871_) );
	AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2869_), .B(_2870_), .C(_2547__bF_buf0), .Y(_2872_) );
	OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf1), .B(_2620__bF_buf4), .C(divider_aOp_abs_16_), .Y(_2873_) );
	NAND3X1 NAND3X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2745_), .B(_2524_), .C(_2769_), .Y(_2874_) );
	AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2873_), .B(_2874_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .Y(_2876_) );
	NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_15_), .B(_1746__bF_buf1), .Y(_2877_) );
	INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_2877_), .Y(_2878_) );
	NAND3X1 NAND3X1_581 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .B(_2874_), .C(_2873_), .Y(_2879_) );
	AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_2879_), .C(_2876_), .Y(_2880_) );
	OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2880_), .C(_2871_), .Y(_2881_) );
	AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_2865_), .C(_2854_), .Y(_2882_) );
	OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_2827_), .B(_2882_), .C(_2816_), .Y(_2883_) );
	NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_2883_), .B(_2742_), .Y(_2884_) );
	AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2884_), .B(_2732_), .C(_1702_), .Y(divider_divuResult_15_) );
	NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_3193_), .Y(_2886_) );
	INVX8 INVX8_27 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .Y(_2887_) );
	NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .B(_2659_), .Y(_2888_) );
	AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2802_), .B(_2801_), .C(_4999__bF_buf6), .Y(_2889_) );
	AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2818_), .B(_2796_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .Y(_2890_) );
	AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2812_), .B(_2806_), .C(_4100__bF_buf5), .Y(_2891_) );
	AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2822_), .B(_2823_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .Y(_2892_) );
	OAI22X1 OAI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_2891_), .B(_2892_), .C(_2889_), .D(_2890_), .Y(_2893_) );
	NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2893_), .B(_2785_), .Y(_2894_) );
	NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(divider_divuResult_16_bF_buf5), .Y(_2895_) );
	OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf0), .B(_2620__bF_buf3), .C(_2225_), .Y(_2897_) );
	NAND3X1 NAND3X1_582 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_2897_), .C(_2895_), .Y(_2898_) );
	OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_2898_), .B(_2872_), .C(_2871_), .Y(_2899_) );
	AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2865_), .B(_2899_), .C(_2854_), .Y(_2900_) );
	NAND3X1 NAND3X1_583 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_2897_), .C(_2895_), .Y(_2901_) );
	NAND3X1 NAND3X1_584 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_2874_), .C(_2873_), .Y(_2902_) );
	NAND3X1 NAND3X1_585 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_2870_), .C(_2869_), .Y(_2903_) );
	INVX1 INVX1_604 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .Y(_2904_) );
	NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .B(divider_divuResult_16_bF_buf4), .Y(_2905_) );
	INVX1 INVX1_605 ( .gnd(gnd), .vdd(vdd), .A(_2561_), .Y(_2906_) );
	OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_3204__bF_buf4), .B(_2620__bF_buf2), .C(_2906_), .Y(_2908_) );
	NAND3X1 NAND3X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_2908_), .C(_2905_), .Y(_2909_) );
	AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_2901_), .B(_2902_), .C(_2903_), .D(_2909_), .Y(_2910_) );
	NAND3X1 NAND3X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_2910_), .C(_2865_), .Y(_2911_) );
	NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_2911_), .B(_2900_), .Y(_2912_) );
	AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_2894_), .C(_2815_), .Y(_2913_) );
	OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_2913_), .C(_2732_), .Y(_2914_) );
	AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_1757__bF_buf0), .C(_2727_), .Y(_2915_) );
	OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf0), .B(_2915_), .C(_2887__bF_buf4), .Y(_2916_) );
	NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf3), .B(_2914_), .Y(_2917_) );
	NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2917__bF_buf4), .Y(_2919_) );
	NAND3X1 NAND3X1_588 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .B(_2229__bF_buf2), .C(_2919_), .Y(_2920_) );
	AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_2916_), .Y(_2921_) );
	INVX8 INVX8_28 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf1), .Y(_2922_) );
	NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_2622_), .Y(_2923_) );
	INVX1 INVX1_606 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2924_) );
	INVX1 INVX1_607 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .Y(_2925_) );
	OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2856_), .C(_2843_), .Y(_2926_) );
	NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_2926_), .Y(_2927_) );
	NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .B(_2926_), .Y(_2928_) );
	INVX1 INVX1_608 ( .gnd(gnd), .vdd(vdd), .A(_2852_), .Y(_2930_) );
	AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2930_), .B(_2928_), .C(_2927_), .Y(_2931_) );
	AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_2829_), .C(_1735__bF_buf0), .Y(_2932_) );
	AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .B(_2843_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .Y(_2933_) );
	AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_2862_), .C(_2470__bF_buf7), .Y(_2934_) );
	AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2848_), .B(_2851_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .Y(_2935_) );
	OAI22X1 OAI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_2933_), .B(_2932_), .C(_2934_), .D(_2935_), .Y(_2936_) );
	AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2905_), .B(_2908_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .Y(_2937_) );
	NAND3X1 NAND3X1_589 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_2908_), .C(_2905_), .Y(_2938_) );
	AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .B(_2938_), .C(_2937_), .Y(_2939_) );
	OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_2936_), .B(_2939_), .C(_2931_), .Y(_2941_) );
	AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_2941_), .C(_2815_), .Y(_2942_) );
	AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_2865_), .B(_2910_), .Y(_2943_) );
	NAND3X1 NAND3X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_2943_), .C(_2894_), .Y(_2944_) );
	AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2942_), .B(_2944_), .C(_2925_), .Y(_2945_) );
	OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .B(_2945_), .C(_2924_), .Y(_2946_) );
	AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2946_), .B(_2726_), .C(_2923_), .Y(_2947_) );
	INVX1 INVX1_609 ( .gnd(gnd), .vdd(vdd), .A(_2923_), .Y(_2948_) );
	INVX1 INVX1_610 ( .gnd(gnd), .vdd(vdd), .A(_2726_), .Y(_2949_) );
	INVX1 INVX1_611 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .Y(_2950_) );
	AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .B(_2911_), .C(_2827_), .Y(_2952_) );
	OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .B(_2952_), .C(_2741_), .Y(_2953_) );
	AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2953_), .B(_2950_), .C(_2658_), .Y(_2954_) );
	NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_2948_), .B(_2949_), .C(_2954_), .Y(_2955_) );
	OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_2955_), .B(_2947_), .C(divider_divuResult_15_bF_buf4), .Y(_2956_) );
	OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_2615_), .B(divider_divuResult_16_bF_buf3), .C(_2628_), .Y(_2957_) );
	OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf3), .B(_2957_), .Y(_2958_) );
	NAND3X1 NAND3X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf3), .B(_2958_), .C(_2956_), .Y(_2959_) );
	OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_2949_), .B(_2954_), .C(_2948_), .Y(_2960_) );
	NAND3X1 NAND3X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2923_), .B(_2726_), .C(_2946_), .Y(_2961_) );
	NAND3X1 NAND3X1_593 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf2), .B(_2960_), .C(_2961_), .Y(_2963_) );
	NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(_2957_), .B(_2917__bF_buf3), .Y(_2964_) );
	NAND3X1 NAND3X1_594 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf0), .B(_2964_), .C(_2963_), .Y(_2965_) );
	NAND3X1 NAND3X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2921_), .B(_2965_), .C(_2959_), .Y(_2966_) );
	NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2646_), .Y(_2967_) );
	INVX1 INVX1_612 ( .gnd(gnd), .vdd(vdd), .A(_2967_), .Y(_2968_) );
	INVX1 INVX1_613 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .Y(_2969_) );
	OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_2723_), .B(_2945_), .C(_2657_), .Y(_2970_) );
	NAND3X1 NAND3X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_2969_), .C(_2970_), .Y(_2971_) );
	AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2652_), .B(_2655_), .C(_2950_), .D(_2953_), .Y(_2972_) );
	OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .B(_2972_), .C(_2967_), .Y(_2974_) );
	NAND3X1 NAND3X1_597 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf1), .B(_2974_), .C(_2971_), .Y(_2975_) );
	OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_2394_), .B(divider_divuResult_16_bF_buf2), .C(_2639_), .Y(_2976_) );
	NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2976_), .B(_2917__bF_buf2), .Y(_2977_) );
	NAND3X1 NAND3X1_598 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf2), .B(_2977_), .C(_2975_), .Y(_2978_) );
	OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .B(_2972_), .C(_2968_), .Y(_2979_) );
	NAND3X1 NAND3X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2967_), .B(_2969_), .C(_2970_), .Y(_2980_) );
	AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_2979_), .C(_2917__bF_buf1), .Y(_2981_) );
	INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(_2977_), .Y(_2982_) );
	OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2981_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .Y(_2983_) );
	INVX1 INVX1_614 ( .gnd(gnd), .vdd(vdd), .A(_2657_), .Y(_2985_) );
	NAND3X1 NAND3X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2985_), .B(_2950_), .C(_2953_), .Y(_2986_) );
	INVX1 INVX1_615 ( .gnd(gnd), .vdd(vdd), .A(_2986_), .Y(_2987_) );
	OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_2972_), .B(_2987_), .C(divider_divuResult_15_bF_buf0), .Y(_2988_) );
	NAND3X1 NAND3X1_601 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_2654_), .C(_2917__bF_buf0), .Y(_2989_) );
	NAND3X1 NAND3X1_602 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf0), .B(_2989_), .C(_2988_), .Y(_2990_) );
	NAND3X1 NAND3X1_603 ( .gnd(gnd), .vdd(vdd), .A(_2649_), .B(_2651_), .C(_2917__bF_buf4), .Y(_2991_) );
	NAND3X1 NAND3X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2970_), .B(_2986_), .C(divider_divuResult_15_bF_buf4), .Y(_2992_) );
	NAND3X1 NAND3X1_605 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .B(_2991_), .C(_2992_), .Y(_2993_) );
	AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_2990_), .B(_2993_), .Y(_2994_) );
	NAND3X1 NAND3X1_606 ( .gnd(gnd), .vdd(vdd), .A(_2978_), .B(_2983_), .C(_2994_), .Y(_2996_) );
	NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .B(_2996_), .Y(_2997_) );
	OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .B(divider_divuResult_16_bF_buf1), .C(_2691_), .Y(_2998_) );
	NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_2917__bF_buf3), .Y(_2999_) );
	INVX1 INVX1_616 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .Y(_3000_) );
	AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2692_), .Y(_3001_) );
	OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .B(_2913_), .C(_2721_), .Y(_3002_) );
	NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_2698_), .B(_3002_), .Y(_3003_) );
	NAND3X1 NAND3X1_607 ( .gnd(gnd), .vdd(vdd), .A(_3000_), .B(_3001_), .C(_3003_), .Y(_3004_) );
	INVX1 INVX1_617 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .Y(_3005_) );
	INVX1 INVX1_618 ( .gnd(gnd), .vdd(vdd), .A(_2698_), .Y(_3007_) );
	INVX1 INVX1_619 ( .gnd(gnd), .vdd(vdd), .A(_2740_), .Y(_3008_) );
	OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .B(_2952_), .C(_3008_), .Y(_3009_) );
	AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_2721_), .C(_3007_), .Y(_3010_) );
	OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .B(_3010_), .C(_3005_), .Y(_3011_) );
	NAND3X1 NAND3X1_608 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf3), .B(_3011_), .C(_3004_), .Y(_3012_) );
	NAND3X1 NAND3X1_609 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf3), .B(_2999_), .C(_3012_), .Y(_3013_) );
	OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf2), .B(_2998_), .Y(_3014_) );
	OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .B(_3010_), .C(_3001_), .Y(_3015_) );
	NAND3X1 NAND3X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3000_), .B(_3005_), .C(_3003_), .Y(_3016_) );
	NAND3X1 NAND3X1_611 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf1), .B(_3015_), .C(_3016_), .Y(_3018_) );
	NAND3X1 NAND3X1_612 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .B(_3014_), .C(_3018_), .Y(_3019_) );
	NAND3X1 NAND3X1_613 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(_2721_), .C(_3009_), .Y(_3020_) );
	INVX1 INVX1_620 ( .gnd(gnd), .vdd(vdd), .A(_3020_), .Y(_3021_) );
	OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_3010_), .B(_3021_), .C(divider_divuResult_15_bF_buf0), .Y(_3022_) );
	NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2917__bF_buf2), .Y(_3023_) );
	NAND3X1 NAND3X1_614 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .B(_3023_), .C(_3022_), .Y(_3024_) );
	NAND3X1 NAND3X1_615 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2693_), .C(_2917__bF_buf1), .Y(_3025_) );
	NAND3X1 NAND3X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_3020_), .C(divider_divuResult_15_bF_buf4), .Y(_3026_) );
	NAND3X1 NAND3X1_617 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf2), .B(_3025_), .C(_3026_), .Y(_3027_) );
	NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(_3027_), .B(_3024_), .Y(_3029_) );
	NAND3X1 NAND3X1_618 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_3019_), .C(_3029_), .Y(_3030_) );
	NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_2709_), .B(_2917__bF_buf0), .Y(_3031_) );
	INVX1 INVX1_621 ( .gnd(gnd), .vdd(vdd), .A(_2720_), .Y(_3032_) );
	NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_2736_), .Y(_3033_) );
	OAI22X1 OAI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_2737_), .B(_2739_), .C(_2815_), .D(_2952_), .Y(_3034_) );
	AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_3032_), .C(_3033_), .Y(_3035_) );
	INVX1 INVX1_622 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .Y(_3036_) );
	NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2737_), .B(_2739_), .Y(_3037_) );
	AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2942_), .B(_2944_), .C(_3037_), .Y(_3038_) );
	NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_2720_), .B(_3036_), .C(_3038_), .Y(_3040_) );
	OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_3035_), .B(_3040_), .C(divider_divuResult_15_bF_buf3), .Y(_3041_) );
	NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_3041_), .Y(_3042_) );
	INVX1 INVX1_623 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .Y(_3043_) );
	NAND3X1 NAND3X1_619 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_2944_), .C(_2942_), .Y(_3044_) );
	NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_3044_), .Y(_3045_) );
	NAND3X1 NAND3X1_620 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf2), .B(_2914_), .C(_3045_), .Y(_3046_) );
	NAND3X1 NAND3X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2717_), .B(_2719_), .C(_2917__bF_buf4), .Y(_3047_) );
	NAND3X1 NAND3X1_622 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf2), .B(_3046_), .C(_3047_), .Y(_3048_) );
	OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .B(_3042_), .C(_3048_), .Y(_3049_) );
	OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf2), .B(_3043_), .C(_3049_), .Y(_3051_) );
	AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_3018_), .B(_3014_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .Y(_3052_) );
	AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_3026_), .B(_3025_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .Y(_3053_) );
	AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3053_), .C(_3052_), .Y(_3054_) );
	OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_3030_), .C(_3054_), .Y(_3055_) );
	NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_2990_), .B(_2978_), .Y(_3056_) );
	NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2983_), .B(_3056_), .Y(_3057_) );
	INVX1 INVX1_624 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .Y(_3058_) );
	AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2963_), .B(_2964_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .Y(_3059_) );
	AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .B(_2920_), .C(_3058_), .Y(_3060_) );
	OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .B(_3057_), .C(_3060_), .Y(_3062_) );
	AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_3055_), .C(_3062_), .Y(_3063_) );
	AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_2766_), .C(_1757__bF_buf1), .D(_2914_), .Y(_3064_) );
	NAND3X1 NAND3X1_623 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf0), .B(_2772_), .C(_2778_), .Y(_3065_) );
	INVX1 INVX1_625 ( .gnd(gnd), .vdd(vdd), .A(_2784_), .Y(_3066_) );
	INVX1 INVX1_626 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .Y(_3067_) );
	OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_2797_), .C(_3067_), .Y(_3068_) );
	AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_2799_), .B(_3068_), .C(_2826_), .D(_2912_), .Y(_3069_) );
	OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_3066_), .B(_3069_), .C(_3065_), .Y(_3070_) );
	NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .B(_3070_), .Y(_3071_) );
	INVX1 INVX1_627 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .Y(_3073_) );
	INVX1 INVX1_628 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .Y(_3074_) );
	AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .B(_2911_), .C(_2893_), .Y(_3075_) );
	OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_3074_), .B(_3075_), .C(_2784_), .Y(_3076_) );
	NAND3X1 NAND3X1_624 ( .gnd(gnd), .vdd(vdd), .A(_3065_), .B(_3073_), .C(_3076_), .Y(_3077_) );
	AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3071_), .B(_3077_), .C(_2917__bF_buf3), .Y(_3078_) );
	OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_3078_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .Y(_3079_) );
	INVX1 INVX1_629 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .Y(_3080_) );
	AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_3076_), .B(_3065_), .C(_3073_), .Y(_3081_) );
	INVX1 INVX1_630 ( .gnd(gnd), .vdd(vdd), .A(_3077_), .Y(_3082_) );
	OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_3081_), .B(_3082_), .C(divider_divuResult_15_bF_buf2), .Y(_3084_) );
	NAND3X1 NAND3X1_625 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf2), .B(_3080_), .C(_3084_), .Y(_3085_) );
	NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3066_), .B(_3069_), .Y(_3086_) );
	AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_3086_), .B(_3076_), .Y(_3087_) );
	NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(_2773_), .B(_2917__bF_buf2), .Y(_3088_) );
	OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_2917__bF_buf1), .B(_3087_), .C(_3088_), .Y(_3089_) );
	OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_3089_), .C(_3085_), .Y(_3090_) );
	NAND3X1 NAND3X1_626 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .B(_3080_), .C(_3084_), .Y(_3091_) );
	OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_3078_), .C(_8971__bF_buf1), .Y(_3092_) );
	NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3076_), .B(_3086_), .Y(_3093_) );
	NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .B(divider_divuResult_15_bF_buf1), .Y(_3095_) );
	NAND3X1 NAND3X1_627 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_3088_), .C(_3095_), .Y(_3096_) );
	NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_3087_), .B(divider_divuResult_15_bF_buf0), .Y(_3097_) );
	NAND3X1 NAND3X1_628 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_2778_), .C(_2917__bF_buf0), .Y(_3098_) );
	NAND3X1 NAND3X1_629 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf2), .B(_3098_), .C(_3097_), .Y(_3099_) );
	AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .B(_3099_), .C(_3091_), .D(_3092_), .Y(_3100_) );
	NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .B(_2917__bF_buf4), .Y(_3101_) );
	NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_2819_), .Y(_3102_) );
	NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(_2825_), .Y(_3103_) );
	INVX1 INVX1_631 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .Y(_3104_) );
	OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_3104_), .B(_2882_), .C(_3067_), .Y(_3106_) );
	XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .B(_3102_), .Y(_3107_) );
	NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_3107_), .B(divider_divuResult_15_bF_buf4), .Y(_3108_) );
	AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3108_), .B(_3101_), .C(_4714__bF_buf6), .Y(_3109_) );
	NAND3X1 NAND3X1_630 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf5), .B(_3101_), .C(_3108_), .Y(_3110_) );
	XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_3104_), .Y(_3111_) );
	INVX1 INVX1_632 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .Y(_3112_) );
	NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_3112_), .B(divider_divuResult_15_bF_buf3), .Y(_3113_) );
	NAND3X1 NAND3X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2806_), .B(_2812_), .C(_2917__bF_buf3), .Y(_3114_) );
	NAND3X1 NAND3X1_632 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_3114_), .C(_3113_), .Y(_3115_) );
	AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .B(_3110_), .C(_3109_), .Y(_3117_) );
	AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3079_), .B(_3090_), .C(_3117_), .D(_3100_), .Y(_3118_) );
	NAND3X1 NAND3X1_633 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(_3101_), .C(_3108_), .Y(_3119_) );
	NAND3X1 NAND3X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2796_), .B(_2818_), .C(_2917__bF_buf2), .Y(_3120_) );
	XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_3106_), .B(_3102_), .Y(_3121_) );
	NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_3121_), .B(divider_divuResult_15_bF_buf2), .Y(_3122_) );
	NAND3X1 NAND3X1_635 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf4), .B(_3120_), .C(_3122_), .Y(_3123_) );
	NAND3X1 NAND3X1_636 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_3114_), .C(_3113_), .Y(_3124_) );
	NAND3X1 NAND3X1_637 ( .gnd(gnd), .vdd(vdd), .A(_2822_), .B(_2823_), .C(_2917__bF_buf1), .Y(_3125_) );
	NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .B(divider_divuResult_15_bF_buf1), .Y(_3126_) );
	NAND3X1 NAND3X1_638 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_3125_), .C(_3126_), .Y(_3128_) );
	AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3123_), .B(_3119_), .C(_3124_), .D(_3128_), .Y(_3129_) );
	AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3129_), .Y(_3130_) );
	NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2917__bF_buf0), .Y(_3131_) );
	NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_2858_), .Y(_3132_) );
	NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .B(_2863_), .Y(_3133_) );
	AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_3133_), .Y(_3134_) );
	OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_2930_), .B(_3134_), .C(_3132_), .Y(_3135_) );
	NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2930_), .B(_3134_), .Y(_3136_) );
	OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .B(_2845_), .C(_3136_), .Y(_3137_) );
	NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_3135_), .B(_3137_), .Y(_3139_) );
	NAND3X1 NAND3X1_639 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf0), .B(_2914_), .C(_3139_), .Y(_3140_) );
	NAND3X1 NAND3X1_640 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .B(_3140_), .C(_3131_), .Y(_3141_) );
	NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(_2917__bF_buf4), .Y(_3142_) );
	XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_3132_), .Y(_3143_) );
	NAND3X1 NAND3X1_641 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf3), .B(_2914_), .C(_3143_), .Y(_3144_) );
	NAND3X1 NAND3X1_642 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf4), .B(_3144_), .C(_3142_), .Y(_3145_) );
	NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_3141_), .B(_3145_), .Y(_3146_) );
	INVX1 INVX1_633 ( .gnd(gnd), .vdd(vdd), .A(_3134_), .Y(_3147_) );
	OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_3133_), .Y(_3148_) );
	NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .B(_3147_), .Y(_3150_) );
	NAND3X1 NAND3X1_643 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf2), .B(_3150_), .C(_2914_), .Y(_3151_) );
	OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_2850_), .B(divider_divuResult_16_bF_buf0), .C(_2861_), .Y(_3152_) );
	INVX1 INVX1_634 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .Y(_3153_) );
	NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_3153_), .B(_2917__bF_buf3), .Y(_3154_) );
	NAND3X1 NAND3X1_644 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf7), .B(_3151_), .C(_3154_), .Y(_3155_) );
	INVX1 INVX1_635 ( .gnd(gnd), .vdd(vdd), .A(_3150_), .Y(_3156_) );
	NAND3X1 NAND3X1_645 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf1), .B(_3156_), .C(_2914_), .Y(_3157_) );
	NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .B(_2917__bF_buf2), .Y(_3158_) );
	NAND3X1 NAND3X1_646 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .B(_3157_), .C(_3158_), .Y(_3159_) );
	NAND3X1 NAND3X1_647 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .B(_3159_), .C(_3146_), .Y(_3161_) );
	NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .B(_2938_), .Y(_3162_) );
	XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_3162_), .Y(_3163_) );
	NAND3X1 NAND3X1_648 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf0), .B(_3163_), .C(_2914_), .Y(_3164_) );
	INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(_3164_), .Y(_3165_) );
	AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2869_), .B(_2870_), .C(_1757__bF_buf3), .D(_2914_), .Y(_3166_) );
	NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .B(_3166_), .C(_3165_), .Y(_3167_) );
	OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_3165_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .Y(_3168_) );
	OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_2524_), .B(_2748_), .C(_2897_), .Y(_3169_) );
	INVX1 INVX1_636 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .Y(_3170_) );
	NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3170_), .B(_2917__bF_buf1), .Y(_3172_) );
	NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .B(_2901_), .Y(_3173_) );
	XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3173_), .B(_2877_), .Y(_3174_) );
	NAND3X1 NAND3X1_649 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf2), .B(_3174_), .C(_2914_), .Y(_3175_) );
	AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3172_), .B(_3175_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .Y(_3176_) );
	AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3176_), .B(_3168_), .C(_3167_), .Y(_3177_) );
	OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(divider_divuResult_15_bF_buf0), .C(_3140_), .Y(_3178_) );
	NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_3178_), .Y(_3179_) );
	INVX1 INVX1_637 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .Y(_3180_) );
	AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_3180_), .C(_3179_), .Y(_3181_) );
	OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3161_), .C(_3181_), .Y(_3183_) );
	NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .B(_3183_), .Y(_3184_) );
	NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .B(_3159_), .Y(_3185_) );
	AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_3141_), .B(_3145_), .C(_3185_), .Y(_3186_) );
	NAND3X1 NAND3X1_650 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(_1757__bF_buf1), .C(_2914_), .Y(_3187_) );
	NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_15_), .B(_3187_), .Y(_3188_) );
	NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_2877_), .B(divider_divuResult_15_bF_buf4), .Y(_3189_) );
	AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_3188_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .Y(_3190_) );
	NAND3X1 NAND3X1_651 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .B(_3188_), .C(_3189_), .Y(_3191_) );
	NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_14_), .B(_1746__bF_buf0), .Y(_3192_) );
	INVX1 INVX1_638 ( .gnd(gnd), .vdd(vdd), .A(_3192_), .Y(_3194_) );
	AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_3191_), .B(_3194_), .C(_3190_), .Y(_3195_) );
	NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_3166_), .C(_3165_), .Y(_3196_) );
	INVX1 INVX1_639 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .Y(_3197_) );
	AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .B(_3164_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .Y(_3198_) );
	AOI21X1 AOI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_3172_), .B(_3175_), .C(_2547__bF_buf6), .Y(_3199_) );
	INVX1 INVX1_640 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .Y(_3200_) );
	NAND3X1 NAND3X1_652 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf0), .B(_3200_), .C(_2914_), .Y(_3201_) );
	NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(_2917__bF_buf0), .Y(_3202_) );
	AOI21X1 AOI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3202_), .B(_3201_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .Y(_3203_) );
	OAI22X1 OAI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .B(_3203_), .C(_3196_), .D(_3198_), .Y(_3205_) );
	NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3205_), .Y(_3206_) );
	NAND3X1 NAND3X1_653 ( .gnd(gnd), .vdd(vdd), .A(_3186_), .B(_3206_), .C(_3130_), .Y(_3207_) );
	NAND3X1 NAND3X1_654 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_3207_), .C(_3184_), .Y(_3208_) );
	NAND3X1 NAND3X1_655 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .B(_3031_), .C(_3041_), .Y(_3209_) );
	NAND3X1 NAND3X1_656 ( .gnd(gnd), .vdd(vdd), .A(_2735_), .B(_2708_), .C(_2917__bF_buf4), .Y(_3210_) );
	OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_2913_), .C(_3032_), .Y(_3211_) );
	NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .B(_3211_), .Y(_3212_) );
	AOI21X1 AOI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_3032_), .C(_3036_), .Y(_3213_) );
	OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3212_), .C(divider_divuResult_15_bF_buf3), .Y(_3214_) );
	NAND3X1 NAND3X1_657 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf1), .B(_3210_), .C(_3214_), .Y(_3216_) );
	NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_3209_), .B(_3216_), .Y(_3217_) );
	NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_2738_), .B(_2917__bF_buf3), .Y(_3218_) );
	AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_3044_), .B(_3034_), .Y(_3219_) );
	NAND3X1 NAND3X1_658 ( .gnd(gnd), .vdd(vdd), .A(_1757__bF_buf3), .B(_2914_), .C(_3219_), .Y(_3220_) );
	NAND3X1 NAND3X1_659 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .B(_3220_), .C(_3218_), .Y(_3221_) );
	AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3221_), .Y(_3222_) );
	NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_3217_), .Y(_3223_) );
	NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .B(_3030_), .Y(_3224_) );
	NAND3X1 NAND3X1_660 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_3224_), .C(_3208_), .Y(_3225_) );
	AOI21X1 AOI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3225_), .B(_3063_), .C(_2886_), .Y(divider_divuResult_14_) );
	INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .Y(_3227_) );
	NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3080_), .B(_3084_), .Y(_3228_) );
	INVX1 INVX1_641 ( .gnd(gnd), .vdd(vdd), .A(_3228_), .Y(_3229_) );
	OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf0), .B(_3229_), .C(_3090_), .Y(_3230_) );
	NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .B(_3099_), .Y(_3231_) );
	NAND3X1 NAND3X1_661 ( .gnd(gnd), .vdd(vdd), .A(_3079_), .B(_3085_), .C(_3231_), .Y(_3232_) );
	OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_2917__bF_buf2), .B(_3121_), .C(_3101_), .Y(_3233_) );
	INVX1 INVX1_642 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .Y(_3234_) );
	OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .B(_3233_), .C(_3115_), .Y(_3235_) );
	OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf3), .B(_3234_), .C(_3235_), .Y(_3237_) );
	OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_3237_), .B(_3232_), .C(_3230_), .Y(_3238_) );
	AOI21X1 AOI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_3183_), .B(_3130_), .C(_3238_), .Y(_3239_) );
	INVX1 INVX1_643 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .Y(_3240_) );
	NAND3X1 NAND3X1_662 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .B(_2977_), .C(_2975_), .Y(_3241_) );
	OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2981_), .C(_1944__bF_buf1), .Y(_3242_) );
	NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .B(_2990_), .Y(_3243_) );
	AOI21X1 AOI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_3242_), .B(_3241_), .C(_3243_), .Y(_3244_) );
	NAND3X1 NAND3X1_663 ( .gnd(gnd), .vdd(vdd), .A(_3240_), .B(_3244_), .C(_3224_), .Y(_3245_) );
	OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_3245_), .C(_3063_), .Y(_3246_) );
	NAND3X1 NAND3X1_664 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_3164_), .C(_3197_), .Y(_3247_) );
	OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_3165_), .C(_2470__bF_buf5), .Y(_3248_) );
	OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(divider_divuResult_15_bF_buf2), .C(_3175_), .Y(_3249_) );
	NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_3249_), .Y(_3250_) );
	NAND3X1 NAND3X1_665 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_3175_), .C(_3172_), .Y(_3251_) );
	AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(_3247_), .C(_3251_), .D(_3250_), .Y(_3252_) );
	NAND3X1 NAND3X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3186_), .B(_3252_), .C(_3130_), .Y(_3253_) );
	NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3253_), .C(_3245_), .Y(_3254_) );
	OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_3254_), .B(_3246_), .C(_3227_), .Y(_3255_) );
	OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf4), .B(_2915_), .C(_3255__bF_buf5), .Y(_3256_) );
	AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_1626_), .B(_1659_), .Y(_3259_) );
	NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1615__bF_buf2), .Y(_3260_) );
	INVX8 INVX8_29 ( .gnd(gnd), .vdd(vdd), .A(_3260_), .Y(_3261_) );
	NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_3259_), .B(_3261__bF_buf3), .Y(_3262_) );
	INVX8 INVX8_30 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf2), .Y(_3263_) );
	OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .B(divider_divuResult_15_bF_buf1), .C(_2229__bF_buf1), .Y(_3264_) );
	INVX1 INVX1_644 ( .gnd(gnd), .vdd(vdd), .A(_3264_), .Y(_3265_) );
	INVX1 INVX1_645 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .Y(_3266_) );
	INVX1 INVX1_646 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .Y(_3267_) );
	OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(_3267_), .C(_3118_), .Y(_3268_) );
	NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_15_), .B(_1746__bF_buf5), .Y(_3270_) );
	NAND3X1 NAND3X1_667 ( .gnd(gnd), .vdd(vdd), .A(_2878_), .B(_3270_), .C(divider_divuResult_15_bF_buf0), .Y(_3271_) );
	INVX1 INVX1_647 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_15_), .Y(_3272_) );
	NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_2917__bF_buf1), .Y(_3273_) );
	NAND3X1 NAND3X1_668 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf2), .B(_3273_), .C(_3271_), .Y(_3274_) );
	AOI21X1 AOI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_3271_), .B(_3273_), .C(_1768__bF_buf1), .Y(_3275_) );
	OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_3192_), .B(_3275_), .C(_3274_), .Y(_3276_) );
	NAND3X1 NAND3X1_669 ( .gnd(gnd), .vdd(vdd), .A(_3252_), .B(_3276_), .C(_3186_), .Y(_3277_) );
	NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_3165_), .Y(_3278_) );
	NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf4), .B(_3278_), .Y(_3279_) );
	AOI21X1 AOI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .B(_3164_), .C(_2470__bF_buf3), .Y(_3281_) );
	NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_3249_), .Y(_3282_) );
	OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_3281_), .B(_3282_), .C(_3279_), .Y(_3283_) );
	OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(divider_divuResult_15_bF_buf4), .C(_3144_), .Y(_3284_) );
	NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf3), .B(_3284_), .Y(_3285_) );
	NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_3284_), .Y(_3286_) );
	OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .B(_3286_), .C(_3285_), .Y(_3287_) );
	AOI21X1 AOI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_3186_), .B(_3283_), .C(_3287_), .Y(_3288_) );
	NAND3X1 NAND3X1_670 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_3277_), .C(_3288_), .Y(_3289_) );
	NAND3X1 NAND3X1_671 ( .gnd(gnd), .vdd(vdd), .A(_3268_), .B(_3224_), .C(_3289_), .Y(_3290_) );
	OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_3266_), .B(_3290_), .C(_3063_), .Y(_3292_) );
	AOI21X1 AOI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_3227_), .C(_3265_), .Y(_3293_) );
	OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf3), .B(_3293_), .C(_3263__bF_buf3), .Y(_3294_) );
	NAND3X1 NAND3X1_672 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf1), .B(_2229__bF_buf0), .C(_3256_), .Y(_3295_) );
	AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_3295_), .B(_3294_), .Y(_3296_) );
	INVX1 INVX1_648 ( .gnd(gnd), .vdd(vdd), .A(_2965_), .Y(_3297_) );
	NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .B(_3297_), .Y(_3298_) );
	INVX1 INVX1_649 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .Y(_3299_) );
	INVX1 INVX1_650 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .Y(_3300_) );
	AOI21X1 AOI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_3207_), .C(_3300_), .Y(_3301_) );
	OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3301_), .C(_3244_), .Y(_3303_) );
	AOI21X1 AOI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .B(_3057_), .C(_3299_), .Y(_3304_) );
	INVX1 INVX1_651 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .Y(_3305_) );
	INVX1 INVX1_652 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .Y(_3306_) );
	AOI21X1 AOI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3290_), .B(_3306_), .C(_2996_), .Y(_3307_) );
	NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3305_), .C(_3307_), .Y(_3308_) );
	OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_3304_), .C(divider_divuResult_14_bF_buf4), .Y(_3309_) );
	OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_2957_), .B(divider_divuResult_15_bF_buf3), .C(_2956_), .Y(_3310_) );
	NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_3310_), .B(_3255__bF_buf4), .Y(_3311_) );
	NAND3X1 NAND3X1_673 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf3), .B(_3311_), .C(_3309_), .Y(_3312_) );
	OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_3305_), .B(_3307_), .C(_3298_), .Y(_3314_) );
	NAND3X1 NAND3X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_3057_), .C(_3303_), .Y(_3315_) );
	NAND3X1 NAND3X1_675 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf3), .B(_3314_), .C(_3315_), .Y(_3316_) );
	INVX1 INVX1_653 ( .gnd(gnd), .vdd(vdd), .A(_3310_), .Y(_3317_) );
	NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_3317_), .B(_3255__bF_buf3), .Y(_3318_) );
	NAND3X1 NAND3X1_676 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf0), .B(_3318_), .C(_3316_), .Y(_3319_) );
	NAND3X1 NAND3X1_677 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .B(_3296_), .C(_3312_), .Y(_3320_) );
	OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_2981_), .B(_2982_), .C(_3255__bF_buf2), .Y(_3321_) );
	NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_3241_), .B(_3242_), .Y(_3322_) );
	INVX1 INVX1_654 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .Y(_3323_) );
	INVX1 INVX1_655 ( .gnd(gnd), .vdd(vdd), .A(_2990_), .Y(_3325_) );
	AOI21X1 AOI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3290_), .B(_3306_), .C(_3243_), .Y(_3326_) );
	OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_3326_), .C(_3323_), .Y(_3327_) );
	OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3301_), .C(_2994_), .Y(_3328_) );
	NAND3X1 NAND3X1_678 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_2990_), .C(_3328_), .Y(_3329_) );
	NAND3X1 NAND3X1_679 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf2), .B(_3327_), .C(_3329_), .Y(_3330_) );
	NAND3X1 NAND3X1_680 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf2), .B(_3321_), .C(_3330_), .Y(_3331_) );
	OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_3326_), .C(_3322_), .Y(_3332_) );
	NAND3X1 NAND3X1_681 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_2990_), .C(_3328_), .Y(_3333_) );
	NAND3X1 NAND3X1_682 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf1), .B(_3332_), .C(_3333_), .Y(_3334_) );
	NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2981_), .Y(_3336_) );
	NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3255__bF_buf1), .Y(_3337_) );
	NAND3X1 NAND3X1_683 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf4), .B(_3337_), .C(_3334_), .Y(_3338_) );
	NAND3X1 NAND3X1_684 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_3306_), .C(_3290_), .Y(_3339_) );
	INVX1 INVX1_656 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .Y(_3340_) );
	OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_3326_), .B(_3340_), .C(divider_divuResult_14_bF_buf0), .Y(_3341_) );
	NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_2986_), .B(_2970_), .Y(_3342_) );
	OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_2917__bF_buf0), .B(_3342_), .C(_2991_), .Y(_3343_) );
	INVX1 INVX1_657 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .Y(_3344_) );
	NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_3344_), .B(_3255__bF_buf0), .Y(_3345_) );
	NAND3X1 NAND3X1_685 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .B(_3345_), .C(_3341_), .Y(_3347_) );
	NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .B(_3255__bF_buf5), .Y(_3348_) );
	NAND3X1 NAND3X1_686 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .B(_3339_), .C(divider_divuResult_14_bF_buf4), .Y(_3349_) );
	NAND3X1 NAND3X1_687 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf0), .B(_3348_), .C(_3349_), .Y(_3350_) );
	NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_3347_), .B(_3350_), .Y(_3351_) );
	NAND3X1 NAND3X1_688 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_3338_), .C(_3351_), .Y(_3352_) );
	NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .B(_3320_), .Y(_3353_) );
	OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(divider_divuResult_15_bF_buf2), .C(_3018_), .Y(_3354_) );
	OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf3), .B(_3354_), .Y(_3355_) );
	AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3013_), .Y(_3356_) );
	INVX1 INVX1_658 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .Y(_3358_) );
	INVX1 INVX1_659 ( .gnd(gnd), .vdd(vdd), .A(_3223_), .Y(_3359_) );
	NAND3X1 NAND3X1_689 ( .gnd(gnd), .vdd(vdd), .A(_3359_), .B(_3268_), .C(_3289_), .Y(_3360_) );
	NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_3360_), .Y(_3361_) );
	NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_3029_), .B(_3361_), .Y(_3362_) );
	NAND3X1 NAND3X1_690 ( .gnd(gnd), .vdd(vdd), .A(_3356_), .B(_3358_), .C(_3362_), .Y(_3363_) );
	INVX1 INVX1_660 ( .gnd(gnd), .vdd(vdd), .A(_3356_), .Y(_3364_) );
	INVX1 INVX1_661 ( .gnd(gnd), .vdd(vdd), .A(_3029_), .Y(_3365_) );
	AOI21X1 AOI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_3360_), .B(_3051_), .C(_3365_), .Y(_3366_) );
	OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .B(_3366_), .C(_3364_), .Y(_3367_) );
	NAND3X1 NAND3X1_691 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf2), .B(_3367_), .C(_3363_), .Y(_3369_) );
	NAND3X1 NAND3X1_692 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf4), .B(_3355_), .C(_3369_), .Y(_3370_) );
	OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .B(_3366_), .C(_3356_), .Y(_3371_) );
	NAND3X1 NAND3X1_693 ( .gnd(gnd), .vdd(vdd), .A(_3364_), .B(_3358_), .C(_3362_), .Y(_3372_) );
	NAND3X1 NAND3X1_694 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf1), .B(_3371_), .C(_3372_), .Y(_3373_) );
	NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .B(_3255__bF_buf4), .Y(_3374_) );
	NAND3X1 NAND3X1_695 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf2), .B(_3374_), .C(_3373_), .Y(_3375_) );
	NAND3X1 NAND3X1_696 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_3051_), .C(_3360_), .Y(_3376_) );
	INVX1 INVX1_662 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .Y(_3377_) );
	OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_3377_), .C(divider_divuResult_14_bF_buf0), .Y(_3378_) );
	NAND3X1 NAND3X1_697 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3026_), .C(_3255__bF_buf3), .Y(_3380_) );
	NAND3X1 NAND3X1_698 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_3380_), .C(_3378_), .Y(_3381_) );
	NAND3X1 NAND3X1_699 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3376_), .C(divider_divuResult_14_bF_buf4), .Y(_3382_) );
	NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_3020_), .B(_3003_), .Y(_3383_) );
	OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_2917__bF_buf4), .B(_3383_), .C(_3025_), .Y(_3384_) );
	NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_3255__bF_buf2), .Y(_3385_) );
	NAND3X1 NAND3X1_700 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf2), .B(_3385_), .C(_3382_), .Y(_3386_) );
	NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3386_), .Y(_3387_) );
	NAND3X1 NAND3X1_701 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3375_), .C(_3387_), .Y(_3388_) );
	NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_3043_), .B(_3255__bF_buf1), .Y(_3389_) );
	NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_3208_), .Y(_3391_) );
	NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3391_), .Y(_3392_) );
	NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_3217_), .B(_3392_), .Y(_3393_) );
	INVX1 INVX1_663 ( .gnd(gnd), .vdd(vdd), .A(_3217_), .Y(_3394_) );
	NAND3X1 NAND3X1_702 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3394_), .C(_3391_), .Y(_3395_) );
	NAND3X1 NAND3X1_703 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf3), .B(_3395_), .C(_3393_), .Y(_3396_) );
	AOI21X1 AOI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3396_), .B(_3389_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .Y(_3397_) );
	NAND3X1 NAND3X1_704 ( .gnd(gnd), .vdd(vdd), .A(_3046_), .B(_3047_), .C(_3255__bF_buf0), .Y(_3398_) );
	XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3208_), .B(_3222_), .Y(_3399_) );
	NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .B(divider_divuResult_14_bF_buf2), .Y(_3400_) );
	AOI21X1 AOI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_3398_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .Y(_3402_) );
	NAND3X1 NAND3X1_705 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .B(_3389_), .C(_3396_), .Y(_3403_) );
	AOI21X1 AOI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3403_), .C(_3397_), .Y(_3404_) );
	AOI21X1 AOI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3374_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf1), .Y(_3405_) );
	AOI21X1 AOI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3385_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .Y(_3406_) );
	AOI21X1 AOI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_3375_), .B(_3406_), .C(_3405_), .Y(_3407_) );
	OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_3404_), .B(_3388_), .C(_3407_), .Y(_3408_) );
	OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(divider_divuResult_14_bF_buf1), .C(_3330_), .Y(_3409_) );
	OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_3344_), .B(divider_divuResult_14_bF_buf0), .C(_3349_), .Y(_3410_) );
	NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf4), .B(_3410_), .Y(_3411_) );
	OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf3), .B(_3409_), .C(_3411_), .Y(_3413_) );
	NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .B(_3413_), .Y(_3414_) );
	OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_3265_), .B(divider_divuResult_14_bF_buf4), .C(_2229__bF_buf4), .Y(_3415_) );
	AOI21X1 AOI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(_3318_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .Y(_3416_) );
	OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf2), .B(_3415_), .C(_3416_), .Y(_3417_) );
	AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_3294_), .Y(_3418_) );
	OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_3414_), .B(_3320_), .C(_3418_), .Y(_3419_) );
	AOI21X1 AOI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .B(_3408_), .C(_3419_), .Y(_3420_) );
	NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .B(_3255__bF_buf5), .Y(_3421_) );
	AOI21X1 AOI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_3048_), .C(_3394_), .Y(_3422_) );
	INVX1 INVX1_664 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .Y(_3423_) );
	OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_3422_), .B(_3423_), .C(divider_divuResult_14_bF_buf3), .Y(_3424_) );
	NAND3X1 NAND3X1_706 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf1), .B(_3421_), .C(_3424_), .Y(_3425_) );
	NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(_3425_), .Y(_3426_) );
	NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_3398_), .B(_3400_), .Y(_3427_) );
	XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .B(_1265__bF_buf0), .Y(_3428_) );
	NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_3428_), .C(_3388_), .Y(_3429_) );
	AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3353_), .Y(_3430_) );
	AOI21X1 AOI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_3227_), .C(_3229_), .Y(_3431_) );
	NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .B(_3089_), .Y(_3432_) );
	NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_3091_), .B(_3092_), .Y(_3434_) );
	NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3205_), .C(_3161_), .Y(_3435_) );
	OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_3183_), .B(_3435_), .C(_3129_), .Y(_3436_) );
	AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .B(_3099_), .C(_3237_), .D(_3436_), .Y(_3437_) );
	OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .B(_3437_), .C(_3434_), .Y(_3438_) );
	INVX1 INVX1_665 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3439_) );
	INVX1 INVX1_666 ( .gnd(gnd), .vdd(vdd), .A(_3434_), .Y(_3440_) );
	AOI21X1 AOI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .B(_3277_), .C(_3267_), .Y(_3441_) );
	OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .B(_3441_), .C(_3231_), .Y(_3442_) );
	NAND3X1 NAND3X1_707 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3440_), .C(_3442_), .Y(_3443_) );
	AOI21X1 AOI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_3438_), .B(_3443_), .C(_3255__bF_buf4), .Y(_3445_) );
	OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .B(_3445_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .Y(_3446_) );
	OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_3078_), .C(_3255__bF_buf3), .Y(_3447_) );
	NAND3X1 NAND3X1_708 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3434_), .C(_3442_), .Y(_3448_) );
	OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .B(_3437_), .C(_3440_), .Y(_3449_) );
	NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .B(_3449_), .Y(_3450_) );
	OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_3255__bF_buf2), .B(_3450_), .C(_3447_), .Y(_3451_) );
	INVX1 INVX1_667 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .Y(_3452_) );
	NAND3X1 NAND3X1_709 ( .gnd(gnd), .vdd(vdd), .A(_3452_), .B(_3237_), .C(_3436_), .Y(_3453_) );
	NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(_3453_), .B(_3442_), .Y(_3454_) );
	NAND3X1 NAND3X1_710 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3292_), .C(_3454_), .Y(_3456_) );
	NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .B(_3255__bF_buf1), .Y(_3457_) );
	NAND3X1 NAND3X1_711 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf6), .B(_3456_), .C(_3457_), .Y(_3458_) );
	OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .B(_3451_), .C(_3458_), .Y(_3459_) );
	NAND3X1 NAND3X1_712 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .B(_3449_), .C(divider_divuResult_14_bF_buf2), .Y(_3460_) );
	NAND3X1 NAND3X1_713 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf1), .B(_3447_), .C(_3460_), .Y(_3461_) );
	NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .B(_3446_), .Y(_3462_) );
	AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .B(_3453_), .Y(_3463_) );
	NAND3X1 NAND3X1_714 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3292_), .C(_3463_), .Y(_3464_) );
	INVX1 INVX1_668 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .Y(_3465_) );
	NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(_3255__bF_buf0), .Y(_3467_) );
	NAND3X1 NAND3X1_715 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .B(_3464_), .C(_3467_), .Y(_3468_) );
	NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3468_), .Y(_3469_) );
	NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_3462_), .Y(_3470_) );
	NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_3234_), .B(_3255__bF_buf5), .Y(_3471_) );
	INVX1 INVX1_669 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .Y(_3472_) );
	NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_3119_), .B(_3123_), .Y(_3473_) );
	NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3124_), .Y(_3474_) );
	INVX1 INVX1_670 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3475_) );
	AOI21X1 AOI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .B(_3277_), .C(_3475_), .Y(_3476_) );
	OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_3476_), .C(_3473_), .Y(_3478_) );
	INVX1 INVX1_671 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .Y(_3479_) );
	OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_3183_), .B(_3435_), .C(_3474_), .Y(_3480_) );
	NAND3X1 NAND3X1_716 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .B(_3479_), .C(_3480_), .Y(_3481_) );
	AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_3478_), .B(_3481_), .Y(_3482_) );
	NAND3X1 NAND3X1_717 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3292_), .C(_3482_), .Y(_3483_) );
	NAND3X1 NAND3X1_718 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .B(_3483_), .C(_3471_), .Y(_3484_) );
	INVX1 INVX1_672 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .Y(_3485_) );
	AOI21X1 AOI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3483_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .Y(_3486_) );
	INVX1 INVX1_673 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .Y(_3487_) );
	OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_2917__bF_buf3), .B(_3112_), .C(_3125_), .Y(_3489_) );
	INVX1 INVX1_674 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .Y(_3490_) );
	NAND3X1 NAND3X1_719 ( .gnd(gnd), .vdd(vdd), .A(_3475_), .B(_3277_), .C(_3288_), .Y(_3491_) );
	NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_3491_), .B(_3480_), .Y(_3492_) );
	INVX1 INVX1_675 ( .gnd(gnd), .vdd(vdd), .A(_3492_), .Y(_3493_) );
	NAND3X1 NAND3X1_720 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3493_), .C(_3292_), .Y(_3494_) );
	OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .B(divider_divuResult_14_bF_buf1), .C(_3494_), .Y(_3495_) );
	NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf2), .B(_3495_), .Y(_3496_) );
	AOI21X1 AOI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3487_), .B(_3496_), .C(_3485_), .Y(_3497_) );
	AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3459_), .C(_3497_), .D(_3470_), .Y(_3498_) );
	AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3461_), .Y(_3499_) );
	NAND3X1 NAND3X1_721 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_3456_), .C(_3457_), .Y(_3500_) );
	NAND3X1 NAND3X1_722 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf5), .B(_3464_), .C(_3467_), .Y(_3501_) );
	NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_3500_), .B(_3501_), .Y(_3502_) );
	NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .B(_3255__bF_buf4), .Y(_3503_) );
	NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_3481_), .B(_3478_), .Y(_3504_) );
	NAND3X1 NAND3X1_723 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3292_), .C(_3504_), .Y(_3505_) );
	NAND3X1 NAND3X1_724 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .B(_3505_), .C(_3503_), .Y(_3506_) );
	NAND3X1 NAND3X1_725 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf1), .B(_3483_), .C(_3471_), .Y(_3507_) );
	NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .B(_3495_), .Y(_3508_) );
	NAND3X1 NAND3X1_726 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3492_), .C(_3292_), .Y(_3510_) );
	OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(divider_divuResult_14_bF_buf0), .C(_3510_), .Y(_3511_) );
	NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf1), .B(_3511_), .Y(_3512_) );
	AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_3507_), .C(_3508_), .D(_3512_), .Y(_3513_) );
	NAND3X1 NAND3X1_727 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3513_), .C(_3499_), .Y(_3514_) );
	NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(_3255__bF_buf3), .Y(_3515_) );
	OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .B(divider_divuResult_15_bF_buf1), .C(_3151_), .Y(_3516_) );
	INVX1 INVX1_676 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .Y(_3517_) );
	OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_3283_), .B(_3206_), .C(_3517_), .Y(_3518_) );
	OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .B(_3516_), .C(_3518_), .Y(_3519_) );
	XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_3146_), .Y(_3521_) );
	NAND3X1 NAND3X1_728 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3292_), .C(_3521_), .Y(_3522_) );
	AOI21X1 AOI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3515_), .B(_3522_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .Y(_3523_) );
	INVX1 INVX1_677 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .Y(_3524_) );
	NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_3178_), .B(_3255__bF_buf2), .Y(_3525_) );
	XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_3146_), .Y(_3526_) );
	NAND3X1 NAND3X1_729 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3292_), .C(_3526_), .Y(_3527_) );
	AOI21X1 AOI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3525_), .B(_3527_), .C(_4999__bF_buf3), .Y(_3528_) );
	OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3205_), .C(_3177_), .Y(_3529_) );
	XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3529_), .B(_3185_), .Y(_3530_) );
	INVX1 INVX1_678 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .Y(_3532_) );
	NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(divider_divuResult_14_bF_buf4), .Y(_3533_) );
	NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_3516_), .B(_3255__bF_buf1), .Y(_3534_) );
	NAND3X1 NAND3X1_730 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf1), .B(_3534_), .C(_3533_), .Y(_3535_) );
	OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_3528_), .B(_3535_), .C(_3524_), .Y(_3536_) );
	NAND3X1 NAND3X1_731 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_3527_), .C(_3525_), .Y(_3537_) );
	NAND3X1 NAND3X1_732 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf2), .B(_3522_), .C(_3515_), .Y(_3538_) );
	NAND3X1 NAND3X1_733 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .B(_3534_), .C(_3533_), .Y(_3539_) );
	NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(divider_divuResult_14_bF_buf3), .Y(_3540_) );
	NAND3X1 NAND3X1_734 ( .gnd(gnd), .vdd(vdd), .A(_3151_), .B(_3154_), .C(_3255__bF_buf0), .Y(_3541_) );
	NAND3X1 NAND3X1_735 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf0), .B(_3541_), .C(_3540_), .Y(_3543_) );
	AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .B(_3538_), .C(_3539_), .D(_3543_), .Y(_3544_) );
	NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_3196_), .B(_3198_), .Y(_3545_) );
	NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_3251_), .B(_3250_), .Y(_3546_) );
	AOI21X1 AOI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3276_), .B(_3546_), .C(_3176_), .Y(_3547_) );
	XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .B(_3545_), .Y(_3548_) );
	NAND3X1 NAND3X1_736 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3548_), .C(_3292_), .Y(_3549_) );
	OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3166_), .C(_3255__bF_buf5), .Y(_3550_) );
	NAND3X1 NAND3X1_737 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf6), .B(_3549_), .C(_3550_), .Y(_3551_) );
	AOI21X1 AOI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3550_), .B(_3549_), .C(_1735__bF_buf5), .Y(_3552_) );
	INVX1 INVX1_679 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .Y(_3554_) );
	XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3546_), .Y(_3555_) );
	NAND3X1 NAND3X1_738 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3555_), .C(_3292_), .Y(_3556_) );
	OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_3554_), .B(divider_divuResult_14_bF_buf2), .C(_3556_), .Y(_3557_) );
	NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_3557_), .Y(_3558_) );
	OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_3552_), .B(_3558_), .C(_3551_), .Y(_3559_) );
	AOI21X1 AOI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_3544_), .C(_3536_), .Y(_3560_) );
	OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_3514_), .B(_3560_), .C(_3498_), .Y(_3561_) );
	NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_3190_), .B(_3275_), .Y(_3562_) );
	XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .B(_3192_), .Y(_3563_) );
	INVX1 INVX1_680 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .Y(_3565_) );
	NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .B(divider_divuResult_14_bF_buf1), .Y(_3566_) );
	OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_15_), .B(divider_divuResult_15_bF_buf0), .C(_3271_), .Y(_3567_) );
	NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_3567_), .B(_3255__bF_buf4), .Y(_3568_) );
	NAND3X1 NAND3X1_739 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_3568_), .C(_3566_), .Y(_3569_) );
	INVX1 INVX1_681 ( .gnd(gnd), .vdd(vdd), .A(_3569_), .Y(_3570_) );
	INVX1 INVX1_682 ( .gnd(gnd), .vdd(vdd), .A(_3567_), .Y(_3571_) );
	NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3255__bF_buf3), .Y(_3572_) );
	NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(divider_divuResult_14_bF_buf0), .Y(_3573_) );
	NAND3X1 NAND3X1_740 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .B(_3572_), .C(_3573_), .Y(_3574_) );
	AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_3569_), .B(_3574_), .Y(_3576_) );
	INVX1 INVX1_683 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_14_), .Y(_3577_) );
	NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf0), .B(_3577_), .Y(_3578_) );
	NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_3192_), .B(_3578_), .Y(_3579_) );
	NAND3X1 NAND3X1_741 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3579_), .C(_3292_), .Y(_3580_) );
	NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .B(_3255__bF_buf2), .Y(_3581_) );
	NAND3X1 NAND3X1_742 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf0), .B(_3580_), .C(_3581_), .Y(_3582_) );
	NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_13_), .B(_1746__bF_buf4), .Y(_3583_) );
	AOI21X1 AOI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3581_), .B(_3580_), .C(_1768__bF_buf7), .Y(_3584_) );
	OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_3584_), .C(_3582_), .Y(_3585_) );
	AOI21X1 AOI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_3585_), .B(_3576_), .C(_3570_), .Y(_3587_) );
	INVX1 INVX1_684 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .Y(_3588_) );
	NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(divider_divuResult_14_bF_buf4), .Y(_3589_) );
	NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_3554_), .B(_3255__bF_buf1), .Y(_3590_) );
	NAND3X1 NAND3X1_743 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .B(_3590_), .C(_3589_), .Y(_3591_) );
	NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .B(_3255__bF_buf0), .Y(_3592_) );
	NAND3X1 NAND3X1_744 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_3556_), .C(_3592_), .Y(_3593_) );
	NAND3X1 NAND3X1_745 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .B(_3549_), .C(_3550_), .Y(_3594_) );
	OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(divider_divuResult_14_bF_buf3), .C(_3549_), .Y(_3595_) );
	NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf4), .B(_3595_), .Y(_3596_) );
	AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3591_), .B(_3593_), .C(_3594_), .D(_3596_), .Y(_3598_) );
	NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .B(_3598_), .Y(_3599_) );
	NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3599_), .B(_3514_), .C(_3587_), .Y(_3600_) );
	OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_3561_), .B(_3600_), .C(_3430_), .Y(_3601_) );
	AOI21X1 AOI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_3601_), .B(_3420_), .C(_3262__bF_buf4), .Y(divider_divuResult_13_) );
	OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_3256_), .B(divider_divuResult_13_bF_buf5), .C(_2229__bF_buf3), .Y(_3602_) );
	XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .B(divider_absoluteValue_B_flipSign_result_19_bF_buf2), .Y(_3603_) );
	NAND3X1 NAND3X1_746 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .B(_3311_), .C(_3309_), .Y(_3604_) );
	NAND3X1 NAND3X1_747 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf2), .B(_3318_), .C(_3316_), .Y(_3605_) );
	NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3604_), .Y(_3606_) );
	INVX1 INVX1_685 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .Y(_3608_) );
	INVX1 INVX1_686 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .Y(_3609_) );
	INVX1 INVX1_687 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .Y(_3610_) );
	INVX1 INVX1_688 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3611_) );
	OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf0), .B(_3611_), .C(_3459_), .Y(_3612_) );
	NAND3X1 NAND3X1_748 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3461_), .C(_3502_), .Y(_3613_) );
	NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_3511_), .Y(_3614_) );
	OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .B(_3614_), .C(_3484_), .Y(_3615_) );
	OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_3615_), .B(_3613_), .C(_3612_), .Y(_3616_) );
	AOI21X1 AOI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3483_), .C(_7204__bF_buf0), .Y(_3617_) );
	AOI21X1 AOI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3503_), .B(_3505_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .Y(_3619_) );
	NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(_3255__bF_buf5), .Y(_3620_) );
	AOI21X1 AOI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_3620_), .B(_3494_), .C(_4714__bF_buf0), .Y(_3621_) );
	NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .B(_3255__bF_buf4), .Y(_3622_) );
	AOI21X1 AOI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .B(_3510_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .Y(_3623_) );
	OAI22X1 OAI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3619_), .C(_3621_), .D(_3623_), .Y(_3624_) );
	NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3469_), .C(_3624_), .Y(_3625_) );
	NAND3X1 NAND3X1_749 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .B(_3522_), .C(_3515_), .Y(_3626_) );
	AOI21X1 AOI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3541_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .Y(_3627_) );
	AOI21X1 AOI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3627_), .B(_3626_), .C(_3523_), .Y(_3628_) );
	AOI21X1 AOI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_3515_), .B(_3522_), .C(_4999__bF_buf1), .Y(_3630_) );
	AOI21X1 AOI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_3525_), .B(_3527_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .Y(_3631_) );
	AOI21X1 AOI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3541_), .C(_4100__bF_buf7), .Y(_3632_) );
	AOI21X1 AOI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3533_), .B(_3534_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .Y(_3633_) );
	OAI22X1 OAI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3630_), .B(_3631_), .C(_3633_), .D(_3632_), .Y(_3634_) );
	NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .B(_3595_), .Y(_3635_) );
	NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_3595_), .Y(_3636_) );
	AOI21X1 AOI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3592_), .B(_3556_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .Y(_3637_) );
	AOI21X1 AOI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_3636_), .B(_3637_), .C(_3635_), .Y(_3638_) );
	OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_3638_), .B(_3634_), .C(_3628_), .Y(_3639_) );
	AOI21X1 AOI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3625_), .B(_3639_), .C(_3616_), .Y(_3641_) );
	INVX1 INVX1_689 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .Y(_3642_) );
	INVX1 INVX1_690 ( .gnd(gnd), .vdd(vdd), .A(_3579_), .Y(_3643_) );
	NAND3X1 NAND3X1_750 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3643_), .C(_3292_), .Y(_3644_) );
	NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_14_), .B(_3255__bF_buf3), .Y(_3645_) );
	AOI21X1 AOI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_3645_), .B(_3644_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .Y(_3646_) );
	INVX1 INVX1_691 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .Y(_3647_) );
	NAND3X1 NAND3X1_751 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_3644_), .C(_3645_), .Y(_3648_) );
	AOI21X1 AOI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3648_), .C(_3646_), .Y(_3649_) );
	OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_3649_), .C(_3569_), .Y(_3650_) );
	AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3544_), .Y(_3652_) );
	NAND3X1 NAND3X1_752 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_3652_), .C(_3625_), .Y(_3653_) );
	AOI21X1 AOI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3653_), .C(_3610_), .Y(_3654_) );
	OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3654_), .C(_3609_), .Y(_3655_) );
	AOI21X1 AOI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .B(_3414_), .C(_3608_), .Y(_3656_) );
	NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_3338_), .Y(_3657_) );
	OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .B(_3657_), .C(_3331_), .Y(_3658_) );
	INVX1 INVX1_692 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .Y(_3659_) );
	OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3561_), .C(_3429_), .Y(_3660_) );
	AOI21X1 AOI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_3660_), .B(_3659_), .C(_3352_), .Y(_3661_) );
	NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .B(_3658_), .C(_3661_), .Y(_3663_) );
	OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_3656_), .B(_3663_), .C(divider_divuResult_13_bF_buf4), .Y(_3664_) );
	OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_3317_), .B(divider_divuResult_14_bF_buf2), .C(_3309_), .Y(_3665_) );
	NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3353_), .Y(_3666_) );
	INVX1 INVX1_693 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .Y(_3667_) );
	AOI21X1 AOI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_3604_), .B(_3605_), .C(_3667_), .Y(_3668_) );
	OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3667_), .C(_3294_), .Y(_3669_) );
	AOI21X1 AOI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3668_), .C(_3669_), .Y(_3670_) );
	NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_3670_), .B(_3666_), .Y(_3671_) );
	NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_3625_), .Y(_3672_) );
	NAND3X1 NAND3X1_753 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3672_), .C(_3653_), .Y(_3674_) );
	AOI21X1 AOI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3430_), .C(_3671_), .Y(_3675_) );
	OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf4), .C(_3665_), .Y(_3676_) );
	NAND3X1 NAND3X1_754 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf1), .B(_3676_), .C(_3664_), .Y(_3677_) );
	OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3661_), .C(_3606_), .Y(_3678_) );
	NAND3X1 NAND3X1_755 ( .gnd(gnd), .vdd(vdd), .A(_3608_), .B(_3414_), .C(_3655_), .Y(_3679_) );
	NAND3X1 NAND3X1_756 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf3), .B(_3679_), .C(_3678_), .Y(_3680_) );
	OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf2), .B(_3665_), .Y(_3681_) );
	NAND3X1 NAND3X1_757 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf0), .B(_3681_), .C(_3680_), .Y(_3682_) );
	NAND3X1 NAND3X1_758 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3603_), .C(_3677_), .Y(_3683_) );
	OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf2), .B(_3675__bF_buf3), .C(_3409_), .Y(_3685_) );
	INVX1 INVX1_694 ( .gnd(gnd), .vdd(vdd), .A(_3657_), .Y(_3686_) );
	OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3654_), .C(_3351_), .Y(_3687_) );
	NAND3X1 NAND3X1_759 ( .gnd(gnd), .vdd(vdd), .A(_3686_), .B(_3411_), .C(_3687_), .Y(_3688_) );
	INVX1 INVX1_695 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3689_) );
	INVX1 INVX1_696 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .Y(_3690_) );
	AOI21X1 AOI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_3660_), .B(_3659_), .C(_3690_), .Y(_3691_) );
	OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_3689_), .B(_3691_), .C(_3657_), .Y(_3692_) );
	NAND3X1 NAND3X1_760 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf1), .B(_3688_), .C(_3692_), .Y(_3693_) );
	NAND3X1 NAND3X1_761 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf1), .B(_3685_), .C(_3693_), .Y(_3694_) );
	INVX1 INVX1_697 ( .gnd(gnd), .vdd(vdd), .A(_3685_), .Y(_3696_) );
	INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf1), .Y(_3697_) );
	NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .B(_3429_), .Y(_3698_) );
	OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_3599_), .B(_3587_), .C(_3560_), .Y(_3699_) );
	AOI21X1 AOI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3625_), .C(_3616_), .Y(_3700_) );
	OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_3698_), .B(_3700_), .C(_3420_), .Y(_3701_) );
	NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3701_), .Y(_3702_) );
	OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_3689_), .B(_3691_), .C(_3686_), .Y(_3703_) );
	NAND3X1 NAND3X1_762 ( .gnd(gnd), .vdd(vdd), .A(_3657_), .B(_3411_), .C(_3687_), .Y(_3704_) );
	AOI21X1 AOI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3704_), .C(_3702_), .Y(_3705_) );
	OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3705_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .Y(_3707_) );
	NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .B(_3408_), .C(_3654_), .Y(_3708_) );
	OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .B(_3708_), .C(divider_divuResult_13_bF_buf0), .Y(_3709_) );
	NAND3X1 NAND3X1_763 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_3349_), .C(_3702_), .Y(_3710_) );
	NAND3X1 NAND3X1_764 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf1), .B(_3709_), .C(_3710_), .Y(_3711_) );
	OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf0), .B(_3675__bF_buf2), .C(_3410_), .Y(_3712_) );
	NAND3X1 NAND3X1_765 ( .gnd(gnd), .vdd(vdd), .A(_3690_), .B(_3659_), .C(_3660_), .Y(_3713_) );
	NAND3X1 NAND3X1_766 ( .gnd(gnd), .vdd(vdd), .A(_3713_), .B(_3687_), .C(divider_divuResult_13_bF_buf5), .Y(_3714_) );
	NAND3X1 NAND3X1_767 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf2), .B(_3712_), .C(_3714_), .Y(_3715_) );
	AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_3711_), .B(_3715_), .Y(_3716_) );
	NAND3X1 NAND3X1_768 ( .gnd(gnd), .vdd(vdd), .A(_3694_), .B(_3716_), .C(_3707_), .Y(_3718_) );
	NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3718_), .Y(_3719_) );
	OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .B(divider_divuResult_14_bF_buf1), .C(_3369_), .Y(_3720_) );
	OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf4), .B(_3675__bF_buf1), .C(_3720_), .Y(_3721_) );
	NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3375_), .Y(_3722_) );
	INVX1 INVX1_698 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .Y(_3723_) );
	INVX1 INVX1_699 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3724_) );
	INVX1 INVX1_700 ( .gnd(gnd), .vdd(vdd), .A(_3404_), .Y(_3725_) );
	NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_3428_), .Y(_3726_) );
	INVX1 INVX1_701 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .Y(_3727_) );
	AOI21X1 AOI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3653_), .C(_3727_), .Y(_3729_) );
	OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_3729_), .C(_3387_), .Y(_3730_) );
	NAND3X1 NAND3X1_769 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_3724_), .C(_3730_), .Y(_3731_) );
	OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3561_), .C(_3726_), .Y(_3732_) );
	AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3386_), .C(_3404_), .D(_3732_), .Y(_3733_) );
	OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(_3733_), .C(_3722_), .Y(_3734_) );
	NAND3X1 NAND3X1_770 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf4), .B(_3731_), .C(_3734_), .Y(_3735_) );
	NAND3X1 NAND3X1_771 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf3), .B(_3721_), .C(_3735_), .Y(_3736_) );
	OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf3), .B(_3720_), .Y(_3737_) );
	OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(_3733_), .C(_3723_), .Y(_3738_) );
	NAND3X1 NAND3X1_772 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_3724_), .C(_3730_), .Y(_3740_) );
	NAND3X1 NAND3X1_773 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf2), .B(_3740_), .C(_3738_), .Y(_3741_) );
	NAND3X1 NAND3X1_774 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .B(_3737_), .C(_3741_), .Y(_3742_) );
	NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(_3725_), .C(_3729_), .Y(_3743_) );
	OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_3733_), .B(_3743_), .C(divider_divuResult_13_bF_buf1), .Y(_3744_) );
	NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .B(_3362_), .Y(_3745_) );
	OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_3255__bF_buf2), .B(_3745_), .C(_3385_), .Y(_3746_) );
	INVX1 INVX1_702 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .Y(_3747_) );
	OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf0), .C(_3747_), .Y(_3748_) );
	NAND3X1 NAND3X1_775 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf0), .B(_3748_), .C(_3744_), .Y(_3749_) );
	OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf2), .B(_3675__bF_buf4), .C(_3746_), .Y(_3751_) );
	INVX1 INVX1_703 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3752_) );
	NAND3X1 NAND3X1_776 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_3404_), .C(_3732_), .Y(_3753_) );
	NAND3X1 NAND3X1_777 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3753_), .C(divider_divuResult_13_bF_buf0), .Y(_3754_) );
	NAND3X1 NAND3X1_778 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf3), .B(_3751_), .C(_3754_), .Y(_3755_) );
	NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3749_), .Y(_3756_) );
	NAND3X1 NAND3X1_779 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_3736_), .C(_3742_), .Y(_3757_) );
	INVX1 INVX1_704 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .Y(_3758_) );
	AOI21X1 AOI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3653_), .C(_3428_), .Y(_3759_) );
	OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3759_), .C(_3758_), .Y(_3760_) );
	INVX1 INVX1_705 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .Y(_3762_) );
	INVX1 INVX1_706 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .Y(_3763_) );
	OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3561_), .C(_3763_), .Y(_3764_) );
	NAND3X1 NAND3X1_780 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_3426_), .C(_3764_), .Y(_3765_) );
	NAND3X1 NAND3X1_781 ( .gnd(gnd), .vdd(vdd), .A(_3760_), .B(_3765_), .C(divider_divuResult_13_bF_buf5), .Y(_3766_) );
	NAND3X1 NAND3X1_782 ( .gnd(gnd), .vdd(vdd), .A(_3421_), .B(_3424_), .C(_3702_), .Y(_3767_) );
	NAND3X1 NAND3X1_783 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .B(_3766_), .C(_3767_), .Y(_3768_) );
	AOI21X1 AOI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(_3766_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .Y(_3769_) );
	NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .B(_3700_), .Y(_3770_) );
	NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_3764_), .B(_3770_), .Y(_3771_) );
	NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(divider_divuResult_13_bF_buf4), .Y(_3773_) );
	INVX1 INVX1_707 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .Y(_3774_) );
	OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf1), .B(_3675__bF_buf3), .C(_3774_), .Y(_3775_) );
	NAND3X1 NAND3X1_784 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf0), .B(_3775_), .C(_3773_), .Y(_3776_) );
	INVX1 INVX1_708 ( .gnd(gnd), .vdd(vdd), .A(_3776_), .Y(_3777_) );
	OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_3769_), .B(_3777_), .C(_3768_), .Y(_3778_) );
	AOI21X1 AOI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_3741_), .B(_3737_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .Y(_3779_) );
	AOI21X1 AOI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_3754_), .B(_3751_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .Y(_3780_) );
	AOI21X1 AOI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_3742_), .B(_3780_), .C(_3779_), .Y(_3781_) );
	OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_3778_), .B(_3757_), .C(_3781_), .Y(_3782_) );
	NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_3685_), .B(_3693_), .Y(_3784_) );
	INVX1 INVX1_709 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .Y(_3785_) );
	OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_3410_), .B(divider_divuResult_13_bF_buf3), .C(_3709_), .Y(_3786_) );
	OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf1), .B(_3786_), .C(_3694_), .Y(_3787_) );
	OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf0), .B(_3785_), .C(_3787_), .Y(_3788_) );
	INVX8 INVX8_31 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf1), .Y(_3789_) );
	NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf4), .B(_3602_), .Y(_3790_) );
	INVX1 INVX1_710 ( .gnd(gnd), .vdd(vdd), .A(_3790_), .Y(_3791_) );
	AOI21X1 AOI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_3415_), .C(_2240__bF_buf2), .Y(_3792_) );
	NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf0), .B(_3792_), .Y(_3793_) );
	AOI21X1 AOI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3680_), .B(_3681_), .C(divider_absoluteValue_B_flipSign_result_18_bF_buf4), .Y(_3795_) );
	AOI21X1 AOI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_3793_), .C(_3791_), .Y(_3796_) );
	OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3788_), .C(_3796_), .Y(_3797_) );
	AOI21X1 AOI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .B(_3782_), .C(_3797_), .Y(_3798_) );
	NAND3X1 NAND3X1_785 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .B(_3721_), .C(_3735_), .Y(_3799_) );
	NAND3X1 NAND3X1_786 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf2), .B(_3737_), .C(_3741_), .Y(_3800_) );
	NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_3799_), .B(_3800_), .Y(_3801_) );
	NAND3X1 NAND3X1_787 ( .gnd(gnd), .vdd(vdd), .A(_3389_), .B(_3396_), .C(_3702_), .Y(_3802_) );
	NAND3X1 NAND3X1_788 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_3758_), .C(_3764_), .Y(_3803_) );
	OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3759_), .C(_3426_), .Y(_3804_) );
	NAND3X1 NAND3X1_789 ( .gnd(gnd), .vdd(vdd), .A(_3803_), .B(_3804_), .C(divider_divuResult_13_bF_buf2), .Y(_3806_) );
	NAND3X1 NAND3X1_790 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .B(_3806_), .C(_3802_), .Y(_3807_) );
	NAND3X1 NAND3X1_791 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf1), .B(_3766_), .C(_3767_), .Y(_3808_) );
	OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf0), .B(_3675__bF_buf2), .C(_3427_), .Y(_3809_) );
	XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3428_), .Y(_3810_) );
	NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_3810_), .B(divider_divuResult_13_bF_buf1), .Y(_3811_) );
	NAND3X1 NAND3X1_792 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .B(_3809_), .C(_3811_), .Y(_3812_) );
	NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_3776_), .B(_3812_), .Y(_3813_) );
	AOI21X1 AOI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_3807_), .B(_3808_), .C(_3813_), .Y(_3814_) );
	NAND3X1 NAND3X1_793 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_3814_), .C(_3801_), .Y(_3815_) );
	NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3718_), .C(_3815_), .Y(_3817_) );
	OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf4), .B(_3675__bF_buf1), .C(_3451_), .Y(_3818_) );
	AOI21X1 AOI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .B(_3650_), .C(_3639_), .Y(_3819_) );
	OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .B(_3819_), .C(_3615_), .Y(_3820_) );
	NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3820_), .Y(_3821_) );
	NAND3X1 NAND3X1_794 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3499_), .C(_3821_), .Y(_3822_) );
	AOI21X1 AOI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3513_), .C(_3497_), .Y(_3823_) );
	OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_3823_), .C(_3458_), .Y(_3824_) );
	NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3824_), .Y(_3825_) );
	NAND3X1 NAND3X1_795 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf0), .B(_3822_), .C(_3825_), .Y(_3826_) );
	NAND3X1 NAND3X1_796 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .B(_3818_), .C(_3826_), .Y(_3828_) );
	NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_3499_), .B(_3824_), .Y(_3829_) );
	NAND3X1 NAND3X1_797 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3462_), .C(_3821_), .Y(_3830_) );
	NAND3X1 NAND3X1_798 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf5), .B(_3830_), .C(_3829_), .Y(_3831_) );
	OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf0), .C(_3611_), .Y(_3832_) );
	NAND3X1 NAND3X1_799 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_3832_), .C(_3831_), .Y(_3833_) );
	NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_3823_), .Y(_3834_) );
	NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3820_), .Y(_3835_) );
	OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_3834_), .B(_3835_), .C(divider_divuResult_13_bF_buf4), .Y(_3836_) );
	OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_3465_), .B(divider_divuResult_14_bF_buf0), .C(_3456_), .Y(_3837_) );
	OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf2), .B(_3675__bF_buf4), .C(_3837_), .Y(_3839_) );
	NAND3X1 NAND3X1_800 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .B(_3839_), .C(_3836_), .Y(_3840_) );
	XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3823_), .B(_3502_), .Y(_3841_) );
	NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf3), .B(_3841_), .Y(_3842_) );
	INVX1 INVX1_711 ( .gnd(gnd), .vdd(vdd), .A(_3837_), .Y(_3843_) );
	OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf1), .B(_3675__bF_buf3), .C(_3843_), .Y(_3844_) );
	NAND3X1 NAND3X1_801 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf5), .B(_3844_), .C(_3842_), .Y(_3845_) );
	AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .B(_3845_), .C(_3828_), .D(_3833_), .Y(_3846_) );
	OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .B(divider_divuResult_14_bF_buf4), .C(_3483_), .Y(_3847_) );
	INVX1 INVX1_712 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .Y(_3848_) );
	OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf0), .B(_3675__bF_buf2), .C(_3848_), .Y(_3850_) );
	NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3512_), .Y(_3851_) );
	AOI21X1 AOI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3851_), .C(_3614_), .Y(_3852_) );
	OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3619_), .C(_3852_), .Y(_3853_) );
	NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_3507_), .Y(_3854_) );
	NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_3854_), .B(_3852_), .Y(_3855_) );
	INVX1 INVX1_713 ( .gnd(gnd), .vdd(vdd), .A(_3855_), .Y(_3856_) );
	NAND3X1 NAND3X1_802 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3856_), .C(divider_divuResult_13_bF_buf2), .Y(_3857_) );
	NAND3X1 NAND3X1_803 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .B(_3850_), .C(_3857_), .Y(_3858_) );
	OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf4), .B(_3675__bF_buf1), .C(_3847_), .Y(_3859_) );
	INVX1 INVX1_714 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .Y(_3861_) );
	OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_3855_), .B(_3861_), .C(divider_divuResult_13_bF_buf1), .Y(_3862_) );
	NAND3X1 NAND3X1_804 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf4), .B(_3859_), .C(_3862_), .Y(_3863_) );
	OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_3623_), .C(_3699_), .Y(_3864_) );
	INVX1 INVX1_715 ( .gnd(gnd), .vdd(vdd), .A(_3864_), .Y(_3865_) );
	NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_3851_), .B(_3699_), .Y(_3866_) );
	OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .B(_3866_), .C(divider_divuResult_13_bF_buf0), .Y(_3867_) );
	OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf0), .C(_3511_), .Y(_3868_) );
	NAND3X1 NAND3X1_805 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_3868_), .C(_3867_), .Y(_3869_) );
	OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf2), .B(_3675__bF_buf4), .C(_3495_), .Y(_3870_) );
	NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_3866_), .B(_3865_), .Y(_3872_) );
	NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_3872_), .B(divider_divuResult_13_bF_buf5), .Y(_3873_) );
	NAND3X1 NAND3X1_806 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf5), .B(_3870_), .C(_3873_), .Y(_3874_) );
	AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_3869_), .B(_3874_), .C(_3858_), .D(_3863_), .Y(_3875_) );
	NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_3875_), .B(_3846_), .Y(_3876_) );
	OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_3178_), .B(divider_divuResult_14_bF_buf3), .C(_3522_), .Y(_3877_) );
	INVX1 INVX1_716 ( .gnd(gnd), .vdd(vdd), .A(_3877_), .Y(_3878_) );
	OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf1), .B(_3675__bF_buf3), .C(_3878_), .Y(_3879_) );
	NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .B(_3538_), .Y(_3880_) );
	NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3650_), .Y(_3881_) );
	AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3539_), .B(_3543_), .C(_3638_), .D(_3881_), .Y(_3882_) );
	OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_3627_), .B(_3882_), .C(_3880_), .Y(_3883_) );
	INVX1 INVX1_717 ( .gnd(gnd), .vdd(vdd), .A(_3880_), .Y(_3884_) );
	NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_3539_), .B(_3543_), .Y(_3885_) );
	INVX1 INVX1_718 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .Y(_3886_) );
	OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .B(_3587_), .C(_3638_), .Y(_3887_) );
	NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_3887_), .Y(_3888_) );
	NAND3X1 NAND3X1_807 ( .gnd(gnd), .vdd(vdd), .A(_3535_), .B(_3884_), .C(_3888_), .Y(_3889_) );
	NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_3883_), .B(_3889_), .Y(_3890_) );
	NAND3X1 NAND3X1_808 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3701_), .C(_3890_), .Y(_3891_) );
	NAND3X1 NAND3X1_809 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .B(_3879_), .C(_3891_), .Y(_3893_) );
	OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf0), .B(_3675__bF_buf2), .C(_3877_), .Y(_3894_) );
	NAND3X1 NAND3X1_810 ( .gnd(gnd), .vdd(vdd), .A(_3535_), .B(_3880_), .C(_3888_), .Y(_3895_) );
	OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_3627_), .B(_3882_), .C(_3884_), .Y(_3896_) );
	NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_3896_), .B(_3895_), .Y(_3897_) );
	NAND3X1 NAND3X1_811 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3701_), .C(_3897_), .Y(_3898_) );
	NAND3X1 NAND3X1_812 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf6), .B(_3894_), .C(_3898_), .Y(_3899_) );
	XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3887_), .B(_3885_), .Y(_3900_) );
	NAND3X1 NAND3X1_813 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3900_), .C(_3701_), .Y(_3901_) );
	OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_3255__bF_buf1), .B(_3532_), .C(_3541_), .Y(_3902_) );
	INVX1 INVX1_719 ( .gnd(gnd), .vdd(vdd), .A(_3902_), .Y(_3904_) );
	OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf4), .B(_3675__bF_buf1), .C(_3904_), .Y(_3905_) );
	NAND3X1 NAND3X1_814 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf0), .B(_3901_), .C(_3905_), .Y(_3906_) );
	NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_3887_), .Y(_3907_) );
	NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3882_), .B(_3907_), .Y(_3908_) );
	NAND3X1 NAND3X1_815 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3908_), .C(_3701_), .Y(_3909_) );
	OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf0), .C(_3902_), .Y(_3910_) );
	NAND3X1 NAND3X1_816 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .B(_3909_), .C(_3910_), .Y(_3911_) );
	NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3911_), .Y(_3912_) );
	AOI21X1 AOI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_3893_), .B(_3899_), .C(_3912_), .Y(_3913_) );
	NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(_3591_), .Y(_3915_) );
	AOI21X1 AOI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_3915_), .C(_3637_), .Y(_3916_) );
	NAND3X1 NAND3X1_817 ( .gnd(gnd), .vdd(vdd), .A(_3551_), .B(_3636_), .C(_3916_), .Y(_3917_) );
	INVX1 INVX1_720 ( .gnd(gnd), .vdd(vdd), .A(_3915_), .Y(_3918_) );
	OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_3918_), .B(_3587_), .C(_3558_), .Y(_3919_) );
	OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_3635_), .B(_3552_), .C(_3919_), .Y(_3920_) );
	NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .B(_3920_), .Y(_3921_) );
	INVX1 INVX1_721 ( .gnd(gnd), .vdd(vdd), .A(_3921_), .Y(_3922_) );
	NAND3X1 NAND3X1_818 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3701_), .C(_3922_), .Y(_3923_) );
	OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf2), .B(_3675__bF_buf4), .C(_3595_), .Y(_3924_) );
	NAND3X1 NAND3X1_819 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf6), .B(_3923_), .C(_3924_), .Y(_3926_) );
	AOI21X1 AOI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3924_), .B(_3923_), .C(_4100__bF_buf5), .Y(_3927_) );
	INVX1 INVX1_722 ( .gnd(gnd), .vdd(vdd), .A(_3557_), .Y(_3928_) );
	XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_3918_), .Y(_3929_) );
	NAND3X1 NAND3X1_820 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3929_), .C(_3701_), .Y(_3930_) );
	OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_3928_), .B(divider_divuResult_13_bF_buf4), .C(_3930_), .Y(_3931_) );
	NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_3931_), .Y(_3932_) );
	OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_3927_), .B(_3932_), .C(_3926_), .Y(_3933_) );
	NAND3X1 NAND3X1_821 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf5), .B(_3879_), .C(_3891_), .Y(_3934_) );
	AOI21X1 AOI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_3879_), .C(_4714__bF_buf4), .Y(_3935_) );
	OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3935_), .C(_3934_), .Y(_3937_) );
	AOI21X1 AOI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3933_), .C(_3937_), .Y(_3938_) );
	NAND3X1 NAND3X1_822 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf3), .B(_3850_), .C(_3857_), .Y(_3939_) );
	AOI21X1 AOI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_3857_), .B(_3850_), .C(_8971__bF_buf2), .Y(_3940_) );
	NAND3X1 NAND3X1_823 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf4), .B(_3868_), .C(_3867_), .Y(_3941_) );
	AOI21X1 AOI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_3939_), .B(_3941_), .C(_3940_), .Y(_3942_) );
	NAND3X1 NAND3X1_824 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf4), .B(_3818_), .C(_3826_), .Y(_3943_) );
	AOI21X1 AOI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_3826_), .B(_3818_), .C(_1265__bF_buf3), .Y(_3944_) );
	NAND3X1 NAND3X1_825 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf4), .B(_3839_), .C(_3836_), .Y(_3945_) );
	OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_3945_), .B(_3944_), .C(_3943_), .Y(_3946_) );
	AOI21X1 AOI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_3846_), .B(_3942_), .C(_3946_), .Y(_3948_) );
	OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_3876_), .B(_3938_), .C(_3948_), .Y(_3949_) );
	OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_3255__bF_buf0), .B(_3565_), .C(_3572_), .Y(_3950_) );
	XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3576_), .B(_3649_), .Y(_3951_) );
	INVX1 INVX1_723 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .Y(_3952_) );
	NAND3X1 NAND3X1_826 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3952_), .C(_3701_), .Y(_3953_) );
	OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(divider_divuResult_13_bF_buf3), .C(_3953_), .Y(_3954_) );
	NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_3954_), .Y(_3955_) );
	NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .B(_3584_), .Y(_3956_) );
	XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3956_), .B(_3583_), .Y(_3957_) );
	INVX1 INVX1_724 ( .gnd(gnd), .vdd(vdd), .A(_3957_), .Y(_3959_) );
	NAND3X1 NAND3X1_827 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3959_), .C(_3701_), .Y(_3960_) );
	OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_14_), .B(divider_divuResult_14_bF_buf2), .C(_3580_), .Y(_3961_) );
	OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf1), .B(_3675__bF_buf3), .C(_3961_), .Y(_3962_) );
	NAND3X1 NAND3X1_828 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_3960_), .C(_3962_), .Y(_3963_) );
	OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_3255__bF_buf5), .B(_3563_), .C(_3568_), .Y(_3964_) );
	OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf0), .B(_3675__bF_buf2), .C(_3964_), .Y(_3965_) );
	NAND3X1 NAND3X1_829 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_3953_), .C(_3965_), .Y(_3966_) );
	NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_3963_), .B(_3966_), .Y(_3967_) );
	NAND3X1 NAND3X1_830 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .B(_3953_), .C(_3965_), .Y(_3968_) );
	NAND3X1 NAND3X1_831 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3951_), .C(_3701_), .Y(_3970_) );
	OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf4), .B(_3675__bF_buf1), .C(_3950_), .Y(_3971_) );
	NAND3X1 NAND3X1_832 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf7), .B(_3970_), .C(_3971_), .Y(_3972_) );
	NAND3X1 NAND3X1_833 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_3960_), .C(_3962_), .Y(_3973_) );
	NAND3X1 NAND3X1_834 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3957_), .C(_3701_), .Y(_3974_) );
	INVX1 INVX1_725 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .Y(_3975_) );
	OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf0), .C(_3975_), .Y(_3976_) );
	NAND3X1 NAND3X1_835 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_3974_), .C(_3976_), .Y(_3977_) );
	AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_3972_), .C(_3973_), .D(_3977_), .Y(_3978_) );
	INVX1 INVX1_726 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_13_), .Y(_3979_) );
	NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .B(_3979_), .Y(_3981_) );
	NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_3981_), .Y(_3982_) );
	NAND3X1 NAND3X1_836 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3982_), .C(_3701_), .Y(_3983_) );
	OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf2), .B(_3675__bF_buf4), .C(_3979_), .Y(_3984_) );
	AOI21X1 AOI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_3984_), .B(_3983_), .C(_1768__bF_buf6), .Y(_3985_) );
	NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_12_), .B(_1746__bF_buf3), .Y(_3986_) );
	NAND3X1 NAND3X1_837 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_3983_), .C(_3984_), .Y(_3987_) );
	AOI21X1 AOI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .B(_3987_), .C(_3985_), .Y(_3988_) );
	AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3955_), .B(_3967_), .C(_3988_), .D(_3978_), .Y(_3989_) );
	NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_3893_), .B(_3899_), .Y(_3990_) );
	AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3911_), .Y(_3992_) );
	NAND3X1 NAND3X1_838 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(_3923_), .C(_3924_), .Y(_3993_) );
	NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf1), .B(_3921_), .C(_3675__bF_buf3), .Y(_3994_) );
	AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3549_), .B(_3550_), .C(_3697_), .D(_3701_), .Y(_3995_) );
	OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_3995_), .B(_3994_), .C(_4100__bF_buf4), .Y(_3996_) );
	INVX1 INVX1_727 ( .gnd(gnd), .vdd(vdd), .A(_3929_), .Y(_3997_) );
	NAND3X1 NAND3X1_839 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3997_), .C(_3701_), .Y(_3998_) );
	OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf0), .B(_3675__bF_buf2), .C(_3928_), .Y(_3999_) );
	NAND3X1 NAND3X1_840 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .B(_3998_), .C(_3999_), .Y(_4000_) );
	OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf4), .B(_3675__bF_buf1), .C(_3557_), .Y(_4001_) );
	NAND3X1 NAND3X1_841 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_3930_), .C(_4001_), .Y(_4003_) );
	AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_4000_), .B(_4003_), .C(_3993_), .D(_3996_), .Y(_4004_) );
	NAND3X1 NAND3X1_842 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .B(_3992_), .C(_4004_), .Y(_4005_) );
	NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_4005_), .C(_3876_), .Y(_4006_) );
	OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .B(_4006_), .C(_3817_), .Y(_4007_) );
	AOI21X1 AOI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_4007_), .B(_3798_), .C(_3182_), .Y(divider_divuResult_12_) );
	INVX8 INVX8_32 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf1), .Y(_4008_) );
	NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_4008__bF_buf5), .Y(_4009_) );
	INVX8 INVX8_33 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .Y(_4010_) );
	INVX8 INVX8_34 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf1), .Y(_4011_) );
	OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_3792_), .B(divider_divuResult_12_bF_buf6), .C(_2229__bF_buf2), .Y(_4013_) );
	NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf3), .B(_4013_), .Y(_4014_) );
	NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_3790_), .B(_3793_), .Y(_4015_) );
	AOI21X1 AOI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3664_), .B(_3676_), .C(_3263__bF_buf0), .Y(_4016_) );
	NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_4015_), .C(_4016_), .Y(_4017_) );
	NAND3X1 NAND3X1_843 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .B(_3685_), .C(_3693_), .Y(_4018_) );
	OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3705_), .C(_2887__bF_buf4), .Y(_4019_) );
	NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3711_), .Y(_4020_) );
	AOI21X1 AOI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_4019_), .B(_4018_), .C(_4020_), .Y(_4021_) );
	NAND3X1 NAND3X1_844 ( .gnd(gnd), .vdd(vdd), .A(_4017_), .B(_4021_), .C(_3782_), .Y(_4022_) );
	AOI21X1 AOI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_3685_), .C(_2887__bF_buf3), .Y(_4024_) );
	AOI21X1 AOI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3694_), .B(_3711_), .C(_4024_), .Y(_4025_) );
	INVX1 INVX1_728 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .Y(_4026_) );
	AOI21X1 AOI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_4017_), .B(_4025_), .C(_4026_), .Y(_4027_) );
	NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(_4027_), .Y(_4028_) );
	NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_3807_), .B(_3808_), .Y(_4029_) );
	AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .B(_3776_), .Y(_4030_) );
	NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_4030_), .B(_4029_), .Y(_4031_) );
	NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_4031_), .B(_3757_), .Y(_4032_) );
	NAND3X1 NAND3X1_845 ( .gnd(gnd), .vdd(vdd), .A(_4021_), .B(_4017_), .C(_4032_), .Y(_4033_) );
	AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_3846_), .B(_3875_), .Y(_4035_) );
	NAND3X1 NAND3X1_846 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3911_), .C(_3990_), .Y(_4036_) );
	NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_3995_), .B(_3994_), .Y(_4037_) );
	OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_3557_), .B(divider_divuResult_13_bF_buf2), .C(_3998_), .Y(_4038_) );
	OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .B(_4038_), .C(_3926_), .Y(_4039_) );
	OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf3), .B(_4037_), .C(_4039_), .Y(_4040_) );
	INVX1 INVX1_729 ( .gnd(gnd), .vdd(vdd), .A(_3937_), .Y(_4041_) );
	OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_4040_), .B(_4036_), .C(_4041_), .Y(_4042_) );
	AOI21X1 AOI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3831_), .B(_3832_), .C(_1265__bF_buf2), .Y(_4043_) );
	AOI21X1 AOI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3826_), .B(_3818_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .Y(_4044_) );
	NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .B(_3845_), .Y(_4046_) );
	OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_4043_), .B(_4044_), .C(_4046_), .Y(_4047_) );
	AOI21X1 AOI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3862_), .B(_3859_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .Y(_4048_) );
	NAND3X1 NAND3X1_847 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .B(_3859_), .C(_3862_), .Y(_4049_) );
	AOI21X1 AOI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3873_), .B(_3870_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .Y(_4050_) );
	OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_4048_), .C(_4049_), .Y(_4051_) );
	INVX1 INVX1_730 ( .gnd(gnd), .vdd(vdd), .A(_3943_), .Y(_4052_) );
	NAND3X1 NAND3X1_848 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .B(_3832_), .C(_3831_), .Y(_4053_) );
	INVX1 INVX1_731 ( .gnd(gnd), .vdd(vdd), .A(_3945_), .Y(_4054_) );
	AOI21X1 AOI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_4053_), .C(_4052_), .Y(_4055_) );
	OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_4051_), .B(_4047_), .C(_4055_), .Y(_4057_) );
	AOI21X1 AOI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4035_), .C(_4057_), .Y(_4058_) );
	INVX1 INVX1_732 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .Y(_4059_) );
	OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_4059_), .C(_3967_), .Y(_4060_) );
	NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_3988_), .B(_3978_), .Y(_4061_) );
	AOI21X1 AOI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_4060_), .B(_4061_), .C(_4005_), .Y(_4062_) );
	NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_4035_), .B(_4062_), .Y(_4063_) );
	AOI21X1 AOI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4063_), .C(_4033_), .Y(_4064_) );
	OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_4028_), .B(_4064_), .C(_3193_), .Y(_4065_) );
	AOI21X1 AOI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_4065__bF_buf4), .B(_3602_), .C(_2240__bF_buf1), .Y(_4066_) );
	NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf0), .B(_4066_), .Y(_4068_) );
	AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_4068_), .B(_4014_), .Y(_4069_) );
	NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_4016_), .Y(_4070_) );
	INVX1 INVX1_733 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .Y(_4071_) );
	AOI21X1 AOI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4063_), .C(_3815_), .Y(_4072_) );
	OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_4072_), .C(_4021_), .Y(_4073_) );
	AOI21X1 AOI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_4073_), .B(_3788_), .C(_4071_), .Y(_4074_) );
	INVX1 INVX1_734 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .Y(_4075_) );
	OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_3949_), .C(_4032_), .Y(_4076_) );
	AOI21X1 AOI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_4075_), .C(_3718_), .Y(_4077_) );
	NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(_4025_), .C(_4077_), .Y(_4079_) );
	OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_4074_), .B(_4079_), .C(divider_divuResult_12_bF_buf5), .Y(_4080_) );
	OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .B(divider_divuResult_13_bF_buf1), .C(_3680_), .Y(_4081_) );
	OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf4), .B(_4081_), .Y(_4082_) );
	NAND3X1 NAND3X1_849 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf3), .B(_4082_), .C(_4080_), .Y(_4083_) );
	OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_4025_), .B(_4077_), .C(_4070_), .Y(_4084_) );
	NAND3X1 NAND3X1_850 ( .gnd(gnd), .vdd(vdd), .A(_4071_), .B(_3788_), .C(_4073_), .Y(_4085_) );
	NAND3X1 NAND3X1_851 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf3), .B(_4085_), .C(_4084_), .Y(_4086_) );
	NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_4081_), .B(_4065__bF_buf3), .Y(_4087_) );
	NAND3X1 NAND3X1_852 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf4), .B(_4087_), .C(_4086_), .Y(_4088_) );
	NAND3X1 NAND3X1_853 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .B(_4088_), .C(_4083_), .Y(_4090_) );
	OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3705_), .C(_4065__bF_buf2), .Y(_4091_) );
	NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .B(_4019_), .Y(_4092_) );
	INVX1 INVX1_735 ( .gnd(gnd), .vdd(vdd), .A(_4092_), .Y(_4093_) );
	INVX1 INVX1_736 ( .gnd(gnd), .vdd(vdd), .A(_3711_), .Y(_4094_) );
	AOI21X1 AOI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_4075_), .C(_4020_), .Y(_4095_) );
	OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_4094_), .B(_4095_), .C(_4093_), .Y(_4096_) );
	OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_4072_), .C(_3716_), .Y(_4097_) );
	NAND3X1 NAND3X1_854 ( .gnd(gnd), .vdd(vdd), .A(_4092_), .B(_3711_), .C(_4097_), .Y(_4098_) );
	NAND3X1 NAND3X1_855 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf2), .B(_4098_), .C(_4096_), .Y(_4099_) );
	NAND3X1 NAND3X1_856 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf3), .B(_4091_), .C(_4099_), .Y(_4101_) );
	OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_4094_), .B(_4095_), .C(_4092_), .Y(_4102_) );
	NAND3X1 NAND3X1_857 ( .gnd(gnd), .vdd(vdd), .A(_4093_), .B(_3711_), .C(_4097_), .Y(_4103_) );
	NAND3X1 NAND3X1_858 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf1), .B(_4103_), .C(_4102_), .Y(_4104_) );
	NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_3785_), .B(_4065__bF_buf1), .Y(_4105_) );
	NAND3X1 NAND3X1_859 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf3), .B(_4105_), .C(_4104_), .Y(_4106_) );
	NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(_3782_), .C(_4072_), .Y(_4107_) );
	OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_4095_), .B(_4107_), .C(divider_divuResult_12_bF_buf0), .Y(_4108_) );
	NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(_4065__bF_buf0), .Y(_4109_) );
	NAND3X1 NAND3X1_860 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf0), .B(_4109_), .C(_4108_), .Y(_4110_) );
	OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf6), .B(_3786_), .Y(_4112_) );
	NAND3X1 NAND3X1_861 ( .gnd(gnd), .vdd(vdd), .A(_4020_), .B(_4075_), .C(_4076_), .Y(_4113_) );
	NAND3X1 NAND3X1_862 ( .gnd(gnd), .vdd(vdd), .A(_4113_), .B(_4097_), .C(divider_divuResult_12_bF_buf5), .Y(_4114_) );
	NAND3X1 NAND3X1_863 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf2), .B(_4114_), .C(_4112_), .Y(_4115_) );
	NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_4115_), .B(_4110_), .Y(_4116_) );
	NAND3X1 NAND3X1_864 ( .gnd(gnd), .vdd(vdd), .A(_4101_), .B(_4106_), .C(_4116_), .Y(_4117_) );
	NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_4117_), .B(_4090_), .Y(_4118_) );
	OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_3720_), .B(divider_divuResult_13_bF_buf0), .C(_3741_), .Y(_4119_) );
	NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_4119_), .B(_4065__bF_buf4), .Y(_4120_) );
	OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_3949_), .C(_3814_), .Y(_4121_) );
	AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3749_), .B(_3755_), .C(_3778_), .D(_4121_), .Y(_4123_) );
	OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_3780_), .B(_4123_), .C(_3801_), .Y(_4124_) );
	INVX1 INVX1_737 ( .gnd(gnd), .vdd(vdd), .A(_3801_), .Y(_4125_) );
	INVX1 INVX1_738 ( .gnd(gnd), .vdd(vdd), .A(_3780_), .Y(_4126_) );
	INVX1 INVX1_739 ( .gnd(gnd), .vdd(vdd), .A(_3778_), .Y(_4127_) );
	AOI21X1 AOI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4063_), .C(_4031_), .Y(_4128_) );
	OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_4127_), .B(_4128_), .C(_3756_), .Y(_4129_) );
	NAND3X1 NAND3X1_865 ( .gnd(gnd), .vdd(vdd), .A(_4125_), .B(_4126_), .C(_4129_), .Y(_4130_) );
	NAND3X1 NAND3X1_866 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf4), .B(_4124_), .C(_4130_), .Y(_4131_) );
	NAND3X1 NAND3X1_867 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf0), .B(_4120_), .C(_4131_), .Y(_4132_) );
	AOI21X1 AOI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_4131_), .B(_4120_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .Y(_4134_) );
	NAND3X1 NAND3X1_868 ( .gnd(gnd), .vdd(vdd), .A(_3744_), .B(_3748_), .C(_4065__bF_buf3), .Y(_4135_) );
	INVX1 INVX1_740 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .Y(_4136_) );
	NAND3X1 NAND3X1_869 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_3778_), .C(_4121_), .Y(_4137_) );
	NAND3X1 NAND3X1_870 ( .gnd(gnd), .vdd(vdd), .A(_4137_), .B(_4129_), .C(divider_divuResult_12_bF_buf3), .Y(_4138_) );
	AOI21X1 AOI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_4138_), .B(_4135_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .Y(_4139_) );
	OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_4134_), .C(_4132_), .Y(_4140_) );
	OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf2), .B(_4119_), .Y(_4141_) );
	NAND3X1 NAND3X1_871 ( .gnd(gnd), .vdd(vdd), .A(_3801_), .B(_4126_), .C(_4129_), .Y(_4142_) );
	OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_3780_), .B(_4123_), .C(_4125_), .Y(_4143_) );
	NAND3X1 NAND3X1_872 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf1), .B(_4143_), .C(_4142_), .Y(_4145_) );
	NAND3X1 NAND3X1_873 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf0), .B(_4141_), .C(_4145_), .Y(_4146_) );
	NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_4127_), .C(_4128_), .Y(_4147_) );
	OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_4123_), .B(_4147_), .C(divider_divuResult_12_bF_buf0), .Y(_4148_) );
	NAND3X1 NAND3X1_874 ( .gnd(gnd), .vdd(vdd), .A(_3751_), .B(_3754_), .C(_4065__bF_buf2), .Y(_4149_) );
	NAND3X1 NAND3X1_875 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .B(_4149_), .C(_4148_), .Y(_4150_) );
	NAND3X1 NAND3X1_876 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf1), .B(_4135_), .C(_4138_), .Y(_4151_) );
	NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_4151_), .B(_4150_), .Y(_4152_) );
	NAND3X1 NAND3X1_877 ( .gnd(gnd), .vdd(vdd), .A(_4146_), .B(_4132_), .C(_4152_), .Y(_4153_) );
	AOI21X1 AOI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4063_), .C(_3813_), .Y(_4154_) );
	OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .B(_4154_), .C(_4029_), .Y(_4156_) );
	INVX1 INVX1_741 ( .gnd(gnd), .vdd(vdd), .A(_4029_), .Y(_4157_) );
	OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_3949_), .C(_4030_), .Y(_4158_) );
	NAND3X1 NAND3X1_878 ( .gnd(gnd), .vdd(vdd), .A(_3776_), .B(_4157_), .C(_4158_), .Y(_4159_) );
	NAND3X1 NAND3X1_879 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .B(_4156_), .C(divider_divuResult_12_bF_buf6), .Y(_4160_) );
	NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_3765_), .B(_3760_), .Y(_4161_) );
	OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_4161_), .C(_3767_), .Y(_4162_) );
	NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .B(_4065__bF_buf1), .Y(_4163_) );
	NAND3X1 NAND3X1_880 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .B(_4163_), .C(_4160_), .Y(_4164_) );
	AOI21X1 AOI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_4160_), .B(_4163_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .Y(_4165_) );
	NAND3X1 NAND3X1_881 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .B(_3775_), .C(_4065__bF_buf0), .Y(_4167_) );
	NAND3X1 NAND3X1_882 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_4063_), .C(_4058_), .Y(_4168_) );
	NAND3X1 NAND3X1_883 ( .gnd(gnd), .vdd(vdd), .A(_4158_), .B(_4168_), .C(divider_divuResult_12_bF_buf5), .Y(_4169_) );
	AOI21X1 AOI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_4167_), .B(_4169_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .Y(_4170_) );
	OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .B(_4165_), .C(_4164_), .Y(_4171_) );
	OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .B(_4153_), .C(_4140_), .Y(_4172_) );
	NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4118_), .Y(_4173_) );
	INVX1 INVX1_742 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .Y(_4174_) );
	NAND3X1 NAND3X1_884 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf3), .B(_4082_), .C(_4080_), .Y(_4175_) );
	NAND3X1 NAND3X1_885 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf2), .B(_4087_), .C(_4086_), .Y(_4176_) );
	AOI21X1 AOI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_4175_), .B(_4176_), .C(_4174_), .Y(_4178_) );
	INVX1 INVX1_743 ( .gnd(gnd), .vdd(vdd), .A(_4106_), .Y(_4179_) );
	OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(divider_divuResult_12_bF_buf4), .C(_4114_), .Y(_4180_) );
	NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf1), .B(_4180_), .Y(_4181_) );
	AOI21X1 AOI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_4101_), .B(_4181_), .C(_4179_), .Y(_4182_) );
	OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_4083_), .B(_4174_), .C(_4014_), .Y(_4183_) );
	AOI21X1 AOI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .B(_4182_), .C(_4183_), .Y(_4184_) );
	AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_4184_), .Y(_4185_) );
	AOI21X1 AOI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_4160_), .B(_4163_), .C(_1505__bF_buf2), .Y(_4186_) );
	INVX1 INVX1_744 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .Y(_4187_) );
	OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .B(divider_divuResult_12_bF_buf3), .C(_4160_), .Y(_4189_) );
	NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf2), .B(_4189_), .Y(_4190_) );
	AOI21X1 AOI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_4167_), .B(_4169_), .C(_1494__bF_buf0), .Y(_4191_) );
	NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_4169_), .B(_4167_), .Y(_4192_) );
	NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_4192_), .Y(_4193_) );
	OAI22X1 OAI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_4191_), .B(_4193_), .C(_4186_), .D(_4190_), .Y(_4194_) );
	NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_4153_), .B(_4194_), .Y(_4195_) );
	AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_4118_), .B(_4195_), .Y(_4196_) );
	OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_3611_), .B(divider_divuResult_13_bF_buf5), .C(_3826_), .Y(_4197_) );
	NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_4197_), .B(_4065__bF_buf4), .Y(_4198_) );
	NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_3828_), .B(_3833_), .Y(_4200_) );
	INVX1 INVX1_745 ( .gnd(gnd), .vdd(vdd), .A(_3875_), .Y(_4201_) );
	AOI21X1 AOI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_3971_), .B(_3970_), .C(_2470__bF_buf5), .Y(_4202_) );
	AOI21X1 AOI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_3965_), .B(_3953_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .Y(_4203_) );
	AOI21X1 AOI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_3976_), .B(_3974_), .C(_2547__bF_buf0), .Y(_4204_) );
	AOI21X1 AOI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_3962_), .B(_3960_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .Y(_4205_) );
	OAI22X1 OAI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_4202_), .B(_4203_), .C(_4204_), .D(_4205_), .Y(_4206_) );
	INVX1 INVX1_746 ( .gnd(gnd), .vdd(vdd), .A(_3982_), .Y(_4207_) );
	NAND3X1 NAND3X1_886 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_4207_), .C(_3701_), .Y(_4208_) );
	OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_3262__bF_buf3), .B(_3675__bF_buf0), .C(divider_aOp_abs_13_), .Y(_4209_) );
	NAND3X1 NAND3X1_887 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .B(_4208_), .C(_4209_), .Y(_4211_) );
	INVX1 INVX1_747 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .Y(_4212_) );
	AOI21X1 AOI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_4209_), .B(_4208_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .Y(_4213_) );
	OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_4212_), .B(_4213_), .C(_4211_), .Y(_4214_) );
	OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_4214_), .B(_4206_), .C(_4060_), .Y(_4215_) );
	NAND3X1 NAND3X1_888 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_4004_), .C(_4215_), .Y(_4216_) );
	AOI21X1 AOI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4216_), .B(_3938_), .C(_4201_), .Y(_4217_) );
	OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_3942_), .B(_4217_), .C(_4046_), .Y(_4218_) );
	NAND3X1 NAND3X1_889 ( .gnd(gnd), .vdd(vdd), .A(_4200_), .B(_3945_), .C(_4218_), .Y(_4219_) );
	INVX1 INVX1_748 ( .gnd(gnd), .vdd(vdd), .A(_4200_), .Y(_4220_) );
	OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4062_), .C(_3875_), .Y(_4222_) );
	AOI22X1 AOI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .B(_3845_), .C(_4051_), .D(_4222_), .Y(_4223_) );
	OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_4223_), .C(_4220_), .Y(_4224_) );
	NAND3X1 NAND3X1_890 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf2), .B(_4224_), .C(_4219_), .Y(_4225_) );
	NAND3X1 NAND3X1_891 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf4), .B(_4198_), .C(_4225_), .Y(_4226_) );
	INVX1 INVX1_749 ( .gnd(gnd), .vdd(vdd), .A(_4197_), .Y(_4227_) );
	NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(_4227_), .B(_4065__bF_buf3), .Y(_4228_) );
	OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_4223_), .C(_4200_), .Y(_4229_) );
	NAND3X1 NAND3X1_892 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(_3945_), .C(_4218_), .Y(_4230_) );
	NAND3X1 NAND3X1_893 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf1), .B(_4229_), .C(_4230_), .Y(_4231_) );
	NAND3X1 NAND3X1_894 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .B(_4228_), .C(_4231_), .Y(_4233_) );
	AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_4233_), .Y(_4234_) );
	INVX1 INVX1_750 ( .gnd(gnd), .vdd(vdd), .A(_4046_), .Y(_4235_) );
	NAND3X1 NAND3X1_895 ( .gnd(gnd), .vdd(vdd), .A(_4235_), .B(_4051_), .C(_4222_), .Y(_4236_) );
	INVX1 INVX1_751 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .Y(_4237_) );
	OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_4223_), .B(_4237_), .C(divider_divuResult_12_bF_buf0), .Y(_4238_) );
	OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_3702_), .C(_3839_), .Y(_4239_) );
	NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_4239_), .B(_4065__bF_buf2), .Y(_4240_) );
	NAND3X1 NAND3X1_896 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .B(_4240_), .C(_4238_), .Y(_4241_) );
	INVX1 INVX1_752 ( .gnd(gnd), .vdd(vdd), .A(_4239_), .Y(_4242_) );
	NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_4242_), .B(_4065__bF_buf1), .Y(_4244_) );
	NAND3X1 NAND3X1_897 ( .gnd(gnd), .vdd(vdd), .A(_4218_), .B(_4236_), .C(divider_divuResult_12_bF_buf6), .Y(_4245_) );
	NAND3X1 NAND3X1_898 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf1), .B(_4244_), .C(_4245_), .Y(_4246_) );
	NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .B(_4246_), .Y(_4247_) );
	OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_3848_), .B(divider_divuResult_13_bF_buf4), .C(_3862_), .Y(_4248_) );
	INVX1 INVX1_753 ( .gnd(gnd), .vdd(vdd), .A(_4248_), .Y(_4249_) );
	NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_3863_), .B(_3858_), .Y(_4250_) );
	NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_3874_), .B(_3869_), .Y(_4251_) );
	OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4062_), .C(_4251_), .Y(_4252_) );
	NAND3X1 NAND3X1_899 ( .gnd(gnd), .vdd(vdd), .A(_4250_), .B(_3941_), .C(_4252_), .Y(_4253_) );
	INVX1 INVX1_754 ( .gnd(gnd), .vdd(vdd), .A(_4250_), .Y(_4255_) );
	INVX1 INVX1_755 ( .gnd(gnd), .vdd(vdd), .A(_4251_), .Y(_4256_) );
	AOI21X1 AOI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_4216_), .B(_3938_), .C(_4256_), .Y(_4257_) );
	OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_4257_), .C(_4255_), .Y(_4258_) );
	NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_4253_), .B(_4258_), .Y(_4259_) );
	NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf5), .B(_4259_), .Y(_4260_) );
	OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_4249_), .B(divider_divuResult_12_bF_buf4), .C(_4260_), .Y(_4261_) );
	NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .B(_4261_), .Y(_4262_) );
	NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_4248_), .B(_4065__bF_buf0), .Y(_4263_) );
	NAND3X1 NAND3X1_900 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf3), .B(_4263_), .C(_4260_), .Y(_4264_) );
	OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(divider_divuResult_13_bF_buf3), .C(_3873_), .Y(_4266_) );
	INVX1 INVX1_756 ( .gnd(gnd), .vdd(vdd), .A(_4266_), .Y(_4267_) );
	NAND3X1 NAND3X1_901 ( .gnd(gnd), .vdd(vdd), .A(_4256_), .B(_3938_), .C(_4216_), .Y(_4268_) );
	NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_4268_), .B(_4252_), .Y(_4269_) );
	INVX1 INVX1_757 ( .gnd(gnd), .vdd(vdd), .A(_4269_), .Y(_4270_) );
	NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_4270_), .B(divider_divuResult_12_bF_buf3), .Y(_4271_) );
	OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_4267_), .B(divider_divuResult_12_bF_buf2), .C(_4271_), .Y(_4272_) );
	NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .B(_4272_), .Y(_4273_) );
	NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_4266_), .B(_4065__bF_buf4), .Y(_4274_) );
	NAND3X1 NAND3X1_902 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf1), .B(_4271_), .C(_4274_), .Y(_4275_) );
	AOI22X1 AOI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_4273_), .B(_4275_), .C(_4262_), .D(_4264_), .Y(_4277_) );
	NAND3X1 NAND3X1_903 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .B(_4247_), .C(_4277_), .Y(_4278_) );
	OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_3702_), .C(_3879_), .Y(_4279_) );
	NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_4279_), .B(_4065__bF_buf3), .Y(_4280_) );
	INVX1 INVX1_758 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .Y(_4281_) );
	INVX1 INVX1_759 ( .gnd(gnd), .vdd(vdd), .A(_4004_), .Y(_4282_) );
	OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_4282_), .B(_3989_), .C(_4040_), .Y(_4283_) );
	NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_3992_), .B(_4283_), .Y(_4284_) );
	AOI21X1 AOI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .B(_3906_), .C(_4281_), .Y(_4285_) );
	OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_3902_), .B(divider_divuResult_13_bF_buf2), .C(_3901_), .Y(_4286_) );
	OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_4286_), .C(_4284_), .Y(_4288_) );
	NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .B(_4288_), .Y(_4289_) );
	OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_4285_), .B(_4289_), .C(divider_divuResult_12_bF_buf1), .Y(_4290_) );
	NAND3X1 NAND3X1_904 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .B(_4280_), .C(_4290_), .Y(_4291_) );
	INVX1 INVX1_760 ( .gnd(gnd), .vdd(vdd), .A(_4279_), .Y(_4292_) );
	NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_4292_), .B(_4065__bF_buf2), .Y(_4293_) );
	NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(_4288_), .Y(_4294_) );
	AOI21X1 AOI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .B(_3906_), .C(_3990_), .Y(_4295_) );
	OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_4294_), .B(_4295_), .C(divider_divuResult_12_bF_buf0), .Y(_4296_) );
	NAND3X1 NAND3X1_905 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_4293_), .C(_4296_), .Y(_4297_) );
	INVX1 INVX1_761 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .Y(_4299_) );
	NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_3992_), .B(_4283_), .Y(_4300_) );
	OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_4299_), .B(_4300_), .C(divider_divuResult_12_bF_buf6), .Y(_4301_) );
	NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_4286_), .B(_4065__bF_buf1), .Y(_4302_) );
	NAND3X1 NAND3X1_906 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_4302_), .C(_4301_), .Y(_4303_) );
	NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_4300_), .B(_4299_), .Y(_4304_) );
	NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_4304_), .B(divider_divuResult_12_bF_buf5), .Y(_4305_) );
	NAND3X1 NAND3X1_907 ( .gnd(gnd), .vdd(vdd), .A(_3901_), .B(_3905_), .C(_4065__bF_buf0), .Y(_4306_) );
	NAND3X1 NAND3X1_908 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf3), .B(_4305_), .C(_4306_), .Y(_4307_) );
	AOI22X1 AOI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_4291_), .B(_4297_), .C(_4303_), .D(_4307_), .Y(_4308_) );
	NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_4037_), .B(_4065__bF_buf4), .Y(_4310_) );
	NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_3993_), .B(_3996_), .Y(_4311_) );
	NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_4000_), .B(_4003_), .Y(_4312_) );
	INVX1 INVX1_762 ( .gnd(gnd), .vdd(vdd), .A(_4312_), .Y(_4313_) );
	OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_4313_), .B(_3989_), .C(_3932_), .Y(_4314_) );
	XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_4314_), .B(_4311_), .Y(_4315_) );
	INVX1 INVX1_763 ( .gnd(gnd), .vdd(vdd), .A(_4315_), .Y(_4316_) );
	NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_4316_), .B(divider_divuResult_12_bF_buf4), .Y(_4317_) );
	AOI21X1 AOI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_4310_), .B(_4317_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .Y(_4318_) );
	INVX1 INVX1_764 ( .gnd(gnd), .vdd(vdd), .A(_4318_), .Y(_4319_) );
	OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_4065__bF_buf3), .B(_4315_), .C(_4310_), .Y(_4321_) );
	NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_4313_), .B(_3989_), .Y(_4322_) );
	NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_4312_), .B(_4215_), .Y(_4323_) );
	NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_4322_), .B(_4323_), .Y(_4324_) );
	NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_4324_), .B(divider_divuResult_12_bF_buf3), .Y(_4325_) );
	NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_3931_), .B(_4065__bF_buf2), .Y(_4326_) );
	AOI21X1 AOI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_4326_), .B(_4325_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .Y(_4327_) );
	OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf6), .B(_4321_), .C(_4327_), .Y(_4328_) );
	NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_4319_), .B(_4328_), .Y(_4329_) );
	AOI21X1 AOI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_4296_), .B(_4293_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .Y(_4330_) );
	INVX1 INVX1_765 ( .gnd(gnd), .vdd(vdd), .A(_4330_), .Y(_4332_) );
	NAND3X1 NAND3X1_909 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .B(_4293_), .C(_4296_), .Y(_4333_) );
	INVX1 INVX1_766 ( .gnd(gnd), .vdd(vdd), .A(_4333_), .Y(_4334_) );
	OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_4286_), .B(divider_divuResult_12_bF_buf2), .C(_4305_), .Y(_4335_) );
	NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf2), .B(_4335_), .Y(_4336_) );
	OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_4336_), .B(_4334_), .C(_4332_), .Y(_4337_) );
	AOI21X1 AOI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_4329_), .B(_4308_), .C(_4337_), .Y(_4338_) );
	NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_4233_), .Y(_4339_) );
	AOI21X1 AOI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .B(_4246_), .C(_4339_), .Y(_4340_) );
	AOI21X1 AOI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_4260_), .B(_4263_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .Y(_4341_) );
	NAND3X1 NAND3X1_910 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .B(_4263_), .C(_4260_), .Y(_4343_) );
	AOI21X1 AOI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_4274_), .B(_4271_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .Y(_4344_) );
	OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_4344_), .B(_4341_), .C(_4343_), .Y(_4345_) );
	INVX1 INVX1_767 ( .gnd(gnd), .vdd(vdd), .A(_4345_), .Y(_4346_) );
	OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_4242_), .B(divider_divuResult_12_bF_buf1), .C(_4238_), .Y(_4347_) );
	OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .B(_4347_), .C(_4226_), .Y(_4348_) );
	AOI22X1 AOI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_4233_), .B(_4348_), .C(_4346_), .D(_4340_), .Y(_4349_) );
	OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_4278_), .B(_4338_), .C(_4349_), .Y(_4350_) );
	NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(_4065__bF_buf1), .Y(_4351_) );
	NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_3798_), .B(_4007_), .Y(_4352_) );
	NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_3972_), .Y(_4354_) );
	NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_3973_), .B(_3977_), .Y(_4355_) );
	INVX1 INVX1_768 ( .gnd(gnd), .vdd(vdd), .A(_4355_), .Y(_4356_) );
	OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_4214_), .B(_4356_), .C(_3963_), .Y(_4357_) );
	XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_4357_), .B(_4354_), .Y(_4358_) );
	NAND3X1 NAND3X1_911 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(_4358_), .C(_4352_), .Y(_4359_) );
	NAND3X1 NAND3X1_912 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_4359_), .C(_4351_), .Y(_4360_) );
	OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_3975_), .B(divider_divuResult_13_bF_buf1), .C(_3960_), .Y(_4361_) );
	INVX1 INVX1_769 ( .gnd(gnd), .vdd(vdd), .A(_4361_), .Y(_4362_) );
	NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_4362_), .B(_4065__bF_buf0), .Y(_4363_) );
	OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_4204_), .B(_4205_), .C(_3988_), .Y(_4365_) );
	NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_4214_), .B(_4356_), .Y(_4366_) );
	NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_4365_), .B(_4366_), .Y(_4367_) );
	OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_4065__bF_buf4), .B(_4367_), .C(_4363_), .Y(_4368_) );
	NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf4), .B(_4368_), .Y(_4369_) );
	INVX1 INVX1_770 ( .gnd(gnd), .vdd(vdd), .A(_4358_), .Y(_4370_) );
	NAND3X1 NAND3X1_913 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(_4370_), .C(_4352_), .Y(_4371_) );
	NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_4059_), .B(_4065__bF_buf3), .Y(_4372_) );
	NAND3X1 NAND3X1_914 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .B(_4371_), .C(_4372_), .Y(_4373_) );
	NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .B(_4373_), .Y(_4374_) );
	OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_4369_), .B(_4374_), .C(_4360_), .Y(_4376_) );
	NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_4367_), .B(divider_divuResult_12_bF_buf0), .Y(_4377_) );
	NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_4361_), .B(_4065__bF_buf2), .Y(_4378_) );
	NAND3X1 NAND3X1_915 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .B(_4377_), .C(_4378_), .Y(_4379_) );
	NAND3X1 NAND3X1_916 ( .gnd(gnd), .vdd(vdd), .A(_4365_), .B(_4366_), .C(divider_divuResult_12_bF_buf6), .Y(_4380_) );
	NAND3X1 NAND3X1_917 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf3), .B(_4363_), .C(_4380_), .Y(_4381_) );
	AOI21X1 AOI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_4379_), .B(_4381_), .C(_4374_), .Y(_4382_) );
	NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_4211_), .B(_3987_), .Y(_4383_) );
	XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_4383_), .B(_3986_), .Y(_4384_) );
	NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(divider_divuResult_12_bF_buf5), .Y(_4385_) );
	OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_13_), .B(divider_divuResult_13_bF_buf0), .C(_3983_), .Y(_4387_) );
	NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .B(_4065__bF_buf1), .Y(_4388_) );
	NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_4388_), .Y(_4389_) );
	INVX1 INVX1_771 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_12_), .Y(_4390_) );
	NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_4390_), .Y(_4391_) );
	NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .B(_4391_), .Y(_4392_) );
	NAND3X1 NAND3X1_918 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(_4392_), .C(_4352_), .Y(_4393_) );
	NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_4390_), .B(_4065__bF_buf0), .Y(_4394_) );
	NAND3X1 NAND3X1_919 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_4393_), .C(_4394_), .Y(_4395_) );
	NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_12_), .B(_4065__bF_buf4), .Y(_4396_) );
	INVX1 INVX1_772 ( .gnd(gnd), .vdd(vdd), .A(_4392_), .Y(_4398_) );
	NAND3X1 NAND3X1_920 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(_4398_), .C(_4352_), .Y(_4399_) );
	NAND3X1 NAND3X1_921 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .B(_4399_), .C(_4396_), .Y(_4400_) );
	NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_11_), .B(_1746__bF_buf2), .Y(_4401_) );
	INVX1 INVX1_773 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .Y(_4402_) );
	NAND3X1 NAND3X1_922 ( .gnd(gnd), .vdd(vdd), .A(_4402_), .B(_4395_), .C(_4400_), .Y(_4403_) );
	MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(_4387_), .S(divider_divuResult_12_bF_buf4), .Y(_4404_) );
	OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_4390_), .B(divider_divuResult_12_bF_buf3), .C(_4399_), .Y(_4405_) );
	AOI22X1 AOI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_4405_), .C(_2547__bF_buf7), .D(_4404_), .Y(_4406_) );
	AOI22X1 AOI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_4389_), .C(_4403_), .D(_4406_), .Y(_4407_) );
	AOI21X1 AOI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4407_), .B(_4382_), .C(_4376_), .Y(_4409_) );
	OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_3994_), .B(_3995_), .C(_4065__bF_buf3), .Y(_4410_) );
	NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_4315_), .B(divider_divuResult_12_bF_buf2), .Y(_4411_) );
	NAND3X1 NAND3X1_923 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .B(_4411_), .C(_4410_), .Y(_4412_) );
	NAND3X1 NAND3X1_924 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_4317_), .C(_4310_), .Y(_4413_) );
	OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_4322_), .B(_4323_), .C(divider_divuResult_12_bF_buf1), .Y(_4414_) );
	NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .B(_4065__bF_buf2), .Y(_4415_) );
	NAND3X1 NAND3X1_925 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .B(_4415_), .C(_4414_), .Y(_4416_) );
	NAND3X1 NAND3X1_926 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_4325_), .C(_4326_), .Y(_4417_) );
	AOI22X1 AOI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_4412_), .B(_4413_), .C(_4416_), .D(_4417_), .Y(_4418_) );
	AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_4308_), .B(_4418_), .Y(_4420_) );
	NAND3X1 NAND3X1_927 ( .gnd(gnd), .vdd(vdd), .A(_4340_), .B(_4277_), .C(_4420_), .Y(_4421_) );
	NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_4409_), .B(_4421_), .Y(_4422_) );
	OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_4422_), .C(_4196_), .Y(_4423_) );
	AOI21X1 AOI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .B(_4185_), .C(_4010__bF_buf4), .Y(divider_divuResult_11_) );
	INVX8 INVX8_35 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf1), .Y(_4424_) );
	NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_4184_), .B(_4173_), .Y(_4425_) );
	NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_4195_), .B(_4118_), .Y(_4426_) );
	NAND3X1 NAND3X1_928 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf0), .B(_4240_), .C(_4238_), .Y(_4427_) );
	NAND3X1 NAND3X1_929 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .B(_4244_), .C(_4245_), .Y(_4428_) );
	NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_4427_), .B(_4428_), .Y(_4430_) );
	AOI21X1 AOI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_4260_), .B(_4263_), .C(_10678__bF_buf2), .Y(_4431_) );
	NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_4249_), .B(_4065__bF_buf1), .Y(_4432_) );
	AOI21X1 AOI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_4252_), .B(_3941_), .C(_4255_), .Y(_4433_) );
	OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .B(_4267_), .C(_4252_), .Y(_4434_) );
	NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_4250_), .B(_4434_), .Y(_4435_) );
	OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_4433_), .B(_4435_), .C(divider_divuResult_12_bF_buf0), .Y(_4436_) );
	AOI21X1 AOI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_4436_), .B(_4432_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .Y(_4437_) );
	AOI21X1 AOI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_4274_), .B(_4271_), .C(_8971__bF_buf0), .Y(_4438_) );
	NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_4269_), .B(divider_divuResult_12_bF_buf6), .Y(_4439_) );
	NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_4267_), .B(_4065__bF_buf0), .Y(_4441_) );
	AOI21X1 AOI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_4441_), .B(_4439_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .Y(_4442_) );
	OAI22X1 OAI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_4438_), .B(_4442_), .C(_4431_), .D(_4437_), .Y(_4443_) );
	NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_4339_), .C(_4443_), .Y(_4444_) );
	AOI21X1 AOI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_4296_), .B(_4293_), .C(_7204__bF_buf2), .Y(_4445_) );
	AOI21X1 AOI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_4290_), .B(_4280_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .Y(_4446_) );
	AOI21X1 AOI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_4306_), .B(_4305_), .C(_4714__bF_buf1), .Y(_4447_) );
	AOI21X1 AOI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_4301_), .B(_4302_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .Y(_4448_) );
	OAI22X1 OAI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_4446_), .C(_4448_), .D(_4447_), .Y(_4449_) );
	NAND3X1 NAND3X1_930 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_4317_), .C(_4310_), .Y(_4450_) );
	AOI21X1 AOI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .B(_4450_), .C(_4318_), .Y(_4452_) );
	AOI21X1 AOI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4306_), .B(_4305_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .Y(_4453_) );
	AOI21X1 AOI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_4453_), .B(_4333_), .C(_4330_), .Y(_4454_) );
	OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_4452_), .B(_4449_), .C(_4454_), .Y(_4455_) );
	NAND3X1 NAND3X1_931 ( .gnd(gnd), .vdd(vdd), .A(_4226_), .B(_4233_), .C(_4247_), .Y(_4456_) );
	OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_4227_), .B(divider_divuResult_12_bF_buf5), .C(_4225_), .Y(_4457_) );
	INVX1 INVX1_774 ( .gnd(gnd), .vdd(vdd), .A(_4457_), .Y(_4458_) );
	OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf3), .B(_4458_), .C(_4348_), .Y(_4459_) );
	OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_4345_), .B(_4456_), .C(_4459_), .Y(_4460_) );
	AOI21X1 AOI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_4444_), .B(_4455_), .C(_4460_), .Y(_4461_) );
	INVX1 INVX1_775 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .Y(_4463_) );
	OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_4362_), .B(divider_divuResult_12_bF_buf4), .C(_4377_), .Y(_4464_) );
	NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .B(_4464_), .Y(_4465_) );
	AOI21X1 AOI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_4465_), .B(_4373_), .C(_4463_), .Y(_4466_) );
	NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_4379_), .B(_4381_), .Y(_4467_) );
	NAND3X1 NAND3X1_932 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .B(_4373_), .C(_4467_), .Y(_4468_) );
	NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_4389_), .Y(_4469_) );
	INVX1 INVX1_776 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_11_), .Y(_4470_) );
	NAND3X1 NAND3X1_933 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_4393_), .C(_4394_), .Y(_4471_) );
	NAND3X1 NAND3X1_934 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf2), .B(_4399_), .C(_4396_), .Y(_4472_) );
	AOI22X1 AOI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(_4470_), .C(_4471_), .D(_4472_), .Y(_4474_) );
	OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_12_), .B(divider_divuResult_12_bF_buf3), .C(_4393_), .Y(_4475_) );
	NAND3X1 NAND3X1_935 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf6), .B(_4385_), .C(_4388_), .Y(_4476_) );
	OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .B(_4475_), .C(_4476_), .Y(_4477_) );
	OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_4477_), .B(_4474_), .C(_4469_), .Y(_4478_) );
	OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_4468_), .B(_4478_), .C(_4466_), .Y(_4479_) );
	NAND3X1 NAND3X1_936 ( .gnd(gnd), .vdd(vdd), .A(_4444_), .B(_4420_), .C(_4479_), .Y(_4480_) );
	AOI21X1 AOI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_4480_), .B(_4461_), .C(_4426_), .Y(_4481_) );
	OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_4425_), .B(_4481_), .C(_4009_), .Y(_4482_) );
	AOI21X1 AOI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4013_), .C(_2240__bF_buf0), .Y(_4483_) );
	INVX1 INVX1_777 ( .gnd(gnd), .vdd(vdd), .A(_4483_), .Y(_4485_) );
	NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf3), .B(_4485_), .Y(_4486_) );
	NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf0), .B(_4483_), .Y(_4487_) );
	AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_4486_), .B(_4487_), .Y(_4488_) );
	NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_4176_), .B(_4175_), .Y(_4489_) );
	INVX1 INVX1_778 ( .gnd(gnd), .vdd(vdd), .A(_4489_), .Y(_4490_) );
	INVX1 INVX1_779 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .Y(_4491_) );
	INVX1 INVX1_780 ( .gnd(gnd), .vdd(vdd), .A(_4117_), .Y(_4492_) );
	OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_4409_), .B(_4421_), .C(_4461_), .Y(_4493_) );
	AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_4493_), .B(_4195_), .Y(_4494_) );
	OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4494_), .C(_4492_), .Y(_4496_) );
	AOI21X1 AOI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .B(_4491_), .C(_4490_), .Y(_4497_) );
	INVX1 INVX1_781 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .Y(_4498_) );
	OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_4422_), .C(_4195_), .Y(_4499_) );
	AOI21X1 AOI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_4499_), .B(_4498_), .C(_4117_), .Y(_4500_) );
	NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4489_), .B(_4182_), .C(_4500_), .Y(_4501_) );
	OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_4501_), .B(_4497_), .C(divider_divuResult_11_bF_buf5), .Y(_4502_) );
	OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_4081_), .B(divider_divuResult_12_bF_buf2), .C(_4080_), .Y(_4503_) );
	AOI21X1 AOI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_4196_), .B(_4493_), .C(_4425_), .Y(_4504_) );
	OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(_4503_), .Y(_4505_) );
	NAND3X1 NAND3X1_937 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf2), .B(_4505_), .C(_4502_), .Y(_4507_) );
	OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .B(_4500_), .C(_4489_), .Y(_4508_) );
	NAND3X1 NAND3X1_938 ( .gnd(gnd), .vdd(vdd), .A(_4490_), .B(_4491_), .C(_4496_), .Y(_4509_) );
	NAND3X1 NAND3X1_939 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf4), .B(_4508_), .C(_4509_), .Y(_4510_) );
	NAND3X1 NAND3X1_940 ( .gnd(gnd), .vdd(vdd), .A(_4080_), .B(_4082_), .C(_4482_), .Y(_4511_) );
	NAND3X1 NAND3X1_941 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf3), .B(_4511_), .C(_4510_), .Y(_4512_) );
	NAND3X1 NAND3X1_942 ( .gnd(gnd), .vdd(vdd), .A(_4512_), .B(_4507_), .C(_4488_), .Y(_4513_) );
	OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_3785_), .B(divider_divuResult_12_bF_buf1), .C(_4099_), .Y(_4514_) );
	OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf2), .B(_4504__bF_buf3), .C(_4514_), .Y(_4515_) );
	INVX1 INVX1_782 ( .gnd(gnd), .vdd(vdd), .A(_4101_), .Y(_4516_) );
	NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_4179_), .B(_4516_), .Y(_4518_) );
	INVX1 INVX1_783 ( .gnd(gnd), .vdd(vdd), .A(_4518_), .Y(_4519_) );
	INVX1 INVX1_784 ( .gnd(gnd), .vdd(vdd), .A(_4181_), .Y(_4520_) );
	INVX1 INVX1_785 ( .gnd(gnd), .vdd(vdd), .A(_4116_), .Y(_4521_) );
	AOI21X1 AOI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_4499_), .B(_4498_), .C(_4521_), .Y(_4522_) );
	OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_4520_), .B(_4522_), .C(_4519_), .Y(_4523_) );
	OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4494_), .C(_4116_), .Y(_4524_) );
	NAND3X1 NAND3X1_943 ( .gnd(gnd), .vdd(vdd), .A(_4518_), .B(_4181_), .C(_4524_), .Y(_4525_) );
	NAND3X1 NAND3X1_944 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf3), .B(_4523_), .C(_4525_), .Y(_4526_) );
	NAND3X1 NAND3X1_945 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf1), .B(_4515_), .C(_4526_), .Y(_4527_) );
	OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_4520_), .B(_4522_), .C(_4518_), .Y(_4529_) );
	NAND3X1 NAND3X1_946 ( .gnd(gnd), .vdd(vdd), .A(_4519_), .B(_4181_), .C(_4524_), .Y(_4530_) );
	NAND3X1 NAND3X1_947 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf2), .B(_4529_), .C(_4530_), .Y(_4531_) );
	OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf1), .B(_4514_), .Y(_4532_) );
	NAND3X1 NAND3X1_948 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf2), .B(_4532_), .C(_4531_), .Y(_4533_) );
	NAND3X1 NAND3X1_949 ( .gnd(gnd), .vdd(vdd), .A(_4521_), .B(_4498_), .C(_4499_), .Y(_4534_) );
	INVX1 INVX1_786 ( .gnd(gnd), .vdd(vdd), .A(_4534_), .Y(_4535_) );
	OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_4522_), .B(_4535_), .C(divider_divuResult_11_bF_buf0), .Y(_4536_) );
	OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf5), .B(_4180_), .Y(_4537_) );
	NAND3X1 NAND3X1_950 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf2), .B(_4537_), .C(_4536_), .Y(_4538_) );
	OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf1), .B(_4504__bF_buf2), .C(_4180_), .Y(_4540_) );
	NAND3X1 NAND3X1_951 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf4), .B(_4534_), .C(_4524_), .Y(_4541_) );
	NAND3X1 NAND3X1_952 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf2), .B(_4540_), .C(_4541_), .Y(_4542_) );
	AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_4538_), .B(_4542_), .Y(_4543_) );
	NAND3X1 NAND3X1_953 ( .gnd(gnd), .vdd(vdd), .A(_4527_), .B(_4533_), .C(_4543_), .Y(_4544_) );
	NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_4544_), .B(_4513_), .Y(_4545_) );
	OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_4119_), .B(divider_divuResult_12_bF_buf0), .C(_4145_), .Y(_4546_) );
	AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_4132_), .B(_4146_), .Y(_4547_) );
	INVX1 INVX1_787 ( .gnd(gnd), .vdd(vdd), .A(_4152_), .Y(_4548_) );
	INVX1 INVX1_788 ( .gnd(gnd), .vdd(vdd), .A(_4194_), .Y(_4549_) );
	OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_4422_), .C(_4549_), .Y(_4551_) );
	AOI21X1 AOI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_4551_), .B(_4171_), .C(_4548_), .Y(_4552_) );
	OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_4552_), .C(_4547_), .Y(_4553_) );
	INVX1 INVX1_789 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .Y(_4554_) );
	INVX1 INVX1_790 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4555_) );
	INVX1 INVX1_791 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(_4556_) );
	AOI21X1 AOI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_4480_), .B(_4461_), .C(_4194_), .Y(_4557_) );
	OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_4556_), .B(_4557_), .C(_4152_), .Y(_4558_) );
	NAND3X1 NAND3X1_954 ( .gnd(gnd), .vdd(vdd), .A(_4554_), .B(_4555_), .C(_4558_), .Y(_4559_) );
	NAND3X1 NAND3X1_955 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf3), .B(_4559_), .C(_4553_), .Y(_4560_) );
	OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_4546_), .B(divider_divuResult_11_bF_buf2), .C(_4560_), .Y(_4562_) );
	OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf0), .B(_4504__bF_buf1), .C(_4546_), .Y(_4563_) );
	NAND3X1 NAND3X1_956 ( .gnd(gnd), .vdd(vdd), .A(_4554_), .B(_4547_), .C(_4558_), .Y(_4564_) );
	OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_4552_), .C(_4555_), .Y(_4565_) );
	NAND3X1 NAND3X1_957 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf1), .B(_4564_), .C(_4565_), .Y(_4566_) );
	NAND3X1 NAND3X1_958 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf0), .B(_4563_), .C(_4566_), .Y(_4567_) );
	NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_4135_), .B(_4138_), .Y(_4568_) );
	NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_4152_), .B(_4556_), .C(_4557_), .Y(_4569_) );
	OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_4552_), .B(_4569_), .C(divider_divuResult_11_bF_buf0), .Y(_4570_) );
	OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_4568_), .B(divider_divuResult_11_bF_buf5), .C(_4570_), .Y(_4571_) );
	OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf4), .B(_4571_), .C(_4567_), .Y(_4573_) );
	OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf4), .B(_4562_), .C(_4573_), .Y(_4574_) );
	NAND3X1 NAND3X1_959 ( .gnd(gnd), .vdd(vdd), .A(_4141_), .B(_4145_), .C(_4482_), .Y(_4575_) );
	NAND3X1 NAND3X1_960 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .B(_4575_), .C(_4560_), .Y(_4576_) );
	NAND3X1 NAND3X1_961 ( .gnd(gnd), .vdd(vdd), .A(_4135_), .B(_4138_), .C(_4482_), .Y(_4577_) );
	NAND3X1 NAND3X1_962 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf3), .B(_4577_), .C(_4570_), .Y(_4578_) );
	OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf4), .B(_4504__bF_buf0), .C(_4568_), .Y(_4579_) );
	NAND3X1 NAND3X1_963 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .B(_4171_), .C(_4551_), .Y(_4580_) );
	NAND3X1 NAND3X1_964 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_4558_), .C(divider_divuResult_11_bF_buf4), .Y(_4581_) );
	NAND3X1 NAND3X1_965 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf3), .B(_4579_), .C(_4581_), .Y(_4582_) );
	NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_4582_), .B(_4578_), .Y(_4584_) );
	NAND3X1 NAND3X1_966 ( .gnd(gnd), .vdd(vdd), .A(_4584_), .B(_4576_), .C(_4567_), .Y(_4585_) );
	INVX1 INVX1_792 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .Y(_4586_) );
	INVX1 INVX1_793 ( .gnd(gnd), .vdd(vdd), .A(_4164_), .Y(_4587_) );
	NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_4165_), .B(_4587_), .Y(_4588_) );
	NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_4191_), .B(_4193_), .Y(_4589_) );
	INVX1 INVX1_794 ( .gnd(gnd), .vdd(vdd), .A(_4589_), .Y(_4590_) );
	OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_4350_), .B(_4422_), .C(_4590_), .Y(_4591_) );
	NAND3X1 NAND3X1_967 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_4588_), .C(_4591_), .Y(_4592_) );
	INVX1 INVX1_795 ( .gnd(gnd), .vdd(vdd), .A(_4588_), .Y(_4593_) );
	AOI21X1 AOI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_4480_), .B(_4461_), .C(_4589_), .Y(_4595_) );
	OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .B(_4595_), .C(_4593_), .Y(_4596_) );
	NAND3X1 NAND3X1_968 ( .gnd(gnd), .vdd(vdd), .A(_4592_), .B(_4596_), .C(divider_divuResult_11_bF_buf3), .Y(_4597_) );
	OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_4189_), .B(divider_divuResult_11_bF_buf2), .C(_4597_), .Y(_4598_) );
	INVX1 INVX1_796 ( .gnd(gnd), .vdd(vdd), .A(_4598_), .Y(_4599_) );
	NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_4590_), .B(_4493_), .Y(_4600_) );
	OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_4600_), .C(divider_divuResult_11_bF_buf1), .Y(_4601_) );
	NAND3X1 NAND3X1_969 ( .gnd(gnd), .vdd(vdd), .A(_4167_), .B(_4169_), .C(_4482_), .Y(_4602_) );
	NAND3X1 NAND3X1_970 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf1), .B(_4602_), .C(_4601_), .Y(_4603_) );
	OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .B(_4598_), .C(_4603_), .Y(_4604_) );
	OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf0), .B(_4599_), .C(_4604_), .Y(_4606_) );
	OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .B(_4606_), .C(_4574_), .Y(_4607_) );
	AOI21X1 AOI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_4531_), .B(_4532_), .C(divider_absoluteValue_B_flipSign_result_19_bF_buf1), .Y(_4608_) );
	INVX1 INVX1_797 ( .gnd(gnd), .vdd(vdd), .A(_4538_), .Y(_4609_) );
	OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_4609_), .B(_4608_), .C(_4533_), .Y(_4610_) );
	INVX1 INVX1_798 ( .gnd(gnd), .vdd(vdd), .A(_4486_), .Y(_4611_) );
	AOI21X1 AOI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_4510_), .B(_4511_), .C(divider_absoluteValue_B_flipSign_result_20_bF_buf2), .Y(_4612_) );
	OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_4612_), .C(_4487_), .Y(_4613_) );
	OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_4610_), .B(_4513_), .C(_4613_), .Y(_4614_) );
	AOI21X1 AOI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_4545_), .B(_4607_), .C(_4614_), .Y(_4615_) );
	NAND3X1 NAND3X1_971 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf1), .B(_4505_), .C(_4502_), .Y(_4617_) );
	NAND3X1 NAND3X1_972 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf1), .B(_4511_), .C(_4510_), .Y(_4618_) );
	NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_4618_), .B(_4617_), .Y(_4619_) );
	NAND3X1 NAND3X1_973 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf0), .B(_4515_), .C(_4526_), .Y(_4620_) );
	NAND3X1 NAND3X1_974 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf0), .B(_4532_), .C(_4531_), .Y(_4621_) );
	NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_4542_), .B(_4538_), .Y(_4622_) );
	AOI21X1 AOI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4621_), .C(_4622_), .Y(_4623_) );
	NAND3X1 NAND3X1_975 ( .gnd(gnd), .vdd(vdd), .A(_4488_), .B(_4623_), .C(_4619_), .Y(_4624_) );
	INVX1 INVX1_799 ( .gnd(gnd), .vdd(vdd), .A(_4189_), .Y(_4625_) );
	OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(_4625_), .Y(_4626_) );
	NAND3X1 NAND3X1_976 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .B(_4626_), .C(_4597_), .Y(_4628_) );
	INVX1 INVX1_800 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .Y(_4629_) );
	OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf2), .B(_4504__bF_buf3), .C(_4189_), .Y(_4630_) );
	OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .B(_4595_), .C(_4588_), .Y(_4631_) );
	NAND3X1 NAND3X1_977 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_4593_), .C(_4591_), .Y(_4632_) );
	NAND3X1 NAND3X1_978 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_4632_), .C(divider_divuResult_11_bF_buf0), .Y(_4633_) );
	NAND3X1 NAND3X1_979 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf4), .B(_4630_), .C(_4633_), .Y(_4634_) );
	INVX1 INVX1_801 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .Y(_4635_) );
	OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf1), .B(_4504__bF_buf2), .C(_4192_), .Y(_4636_) );
	NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_4600_), .Y(_4637_) );
	NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf5), .B(_4637_), .Y(_4639_) );
	NAND3X1 NAND3X1_980 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf1), .B(_4636_), .C(_4639_), .Y(_4640_) );
	AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_4640_), .B(_4603_), .Y(_4641_) );
	OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_4629_), .B(_4635_), .C(_4641_), .Y(_4642_) );
	OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .B(_4642_), .Y(_4643_) );
	NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_4643_), .B(_4624_), .Y(_4644_) );
	OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf0), .B(_4504__bF_buf1), .C(_4457_), .Y(_4645_) );
	AOI21X1 AOI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_4420_), .C(_4455_), .Y(_4646_) );
	OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_4443_), .B(_4646_), .C(_4345_), .Y(_4647_) );
	NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_4247_), .B(_4647_), .Y(_4648_) );
	NAND3X1 NAND3X1_981 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .B(_4427_), .C(_4648_), .Y(_4650_) );
	INVX1 INVX1_802 ( .gnd(gnd), .vdd(vdd), .A(_4427_), .Y(_4651_) );
	NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_4403_), .B(_4406_), .Y(_4652_) );
	NAND3X1 NAND3X1_982 ( .gnd(gnd), .vdd(vdd), .A(_4469_), .B(_4382_), .C(_4652_), .Y(_4653_) );
	NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .B(_4308_), .Y(_4654_) );
	AOI21X1 AOI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_4653_), .B(_4466_), .C(_4654_), .Y(_4655_) );
	OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_4455_), .B(_4655_), .C(_4277_), .Y(_4656_) );
	AOI22X1 AOI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .B(_4246_), .C(_4345_), .D(_4656_), .Y(_4657_) );
	OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_4657_), .C(_4339_), .Y(_4658_) );
	NAND3X1 NAND3X1_983 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf4), .B(_4658_), .C(_4650_), .Y(_4659_) );
	NAND3X1 NAND3X1_984 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .B(_4645_), .C(_4659_), .Y(_4661_) );
	OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_4657_), .C(_4234_), .Y(_4662_) );
	NAND3X1 NAND3X1_985 ( .gnd(gnd), .vdd(vdd), .A(_4339_), .B(_4427_), .C(_4648_), .Y(_4663_) );
	NAND3X1 NAND3X1_986 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf3), .B(_4662_), .C(_4663_), .Y(_4664_) );
	OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf4), .B(_4504__bF_buf0), .C(_4458_), .Y(_4665_) );
	NAND3X1 NAND3X1_987 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf4), .B(_4665_), .C(_4664_), .Y(_4666_) );
	NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_4247_), .B(_4647_), .Y(_4667_) );
	OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .B(_4667_), .C(divider_divuResult_11_bF_buf2), .Y(_4668_) );
	OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(_4347_), .Y(_4669_) );
	NAND3X1 NAND3X1_988 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .B(_4669_), .C(_4668_), .Y(_4670_) );
	NAND3X1 NAND3X1_989 ( .gnd(gnd), .vdd(vdd), .A(_4430_), .B(_4345_), .C(_4656_), .Y(_4672_) );
	NAND3X1 NAND3X1_990 ( .gnd(gnd), .vdd(vdd), .A(_4648_), .B(_4672_), .C(divider_divuResult_11_bF_buf1), .Y(_4673_) );
	INVX1 INVX1_803 ( .gnd(gnd), .vdd(vdd), .A(_4347_), .Y(_4674_) );
	OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf2), .B(_4504__bF_buf3), .C(_4674_), .Y(_4675_) );
	NAND3X1 NAND3X1_991 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf2), .B(_4675_), .C(_4673_), .Y(_4676_) );
	AOI22X1 AOI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_4670_), .B(_4676_), .C(_4661_), .D(_4666_), .Y(_4677_) );
	OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf0), .B(_4261_), .Y(_4678_) );
	NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_4264_), .B(_4262_), .Y(_4679_) );
	INVX1 INVX1_804 ( .gnd(gnd), .vdd(vdd), .A(_4344_), .Y(_4680_) );
	NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_4275_), .B(_4273_), .Y(_4681_) );
	INVX1 INVX1_805 ( .gnd(gnd), .vdd(vdd), .A(_4681_), .Y(_4683_) );
	OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_4646_), .C(_4680_), .Y(_4684_) );
	AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_4684_), .B(_4679_), .Y(_4685_) );
	NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_4679_), .B(_4684_), .Y(_4686_) );
	OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_4686_), .B(_4685_), .C(divider_divuResult_11_bF_buf5), .Y(_4687_) );
	NAND3X1 NAND3X1_992 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .B(_4687_), .C(_4678_), .Y(_4688_) );
	OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf1), .B(_4504__bF_buf2), .C(_4261_), .Y(_4689_) );
	INVX1 INVX1_806 ( .gnd(gnd), .vdd(vdd), .A(_4679_), .Y(_4690_) );
	NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_4690_), .B(_4684_), .Y(_4691_) );
	AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_4684_), .B(_4690_), .Y(_4692_) );
	OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_4691_), .B(_4692_), .C(divider_divuResult_11_bF_buf4), .Y(_4694_) );
	NAND3X1 NAND3X1_993 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_4689_), .C(_4694_), .Y(_4695_) );
	NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_4646_), .Y(_4696_) );
	OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4409_), .C(_4338_), .Y(_4697_) );
	NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_4681_), .B(_4697_), .Y(_4698_) );
	OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_4696_), .B(_4698_), .C(divider_divuResult_11_bF_buf3), .Y(_4699_) );
	INVX1 INVX1_807 ( .gnd(gnd), .vdd(vdd), .A(_4272_), .Y(_4700_) );
	OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf0), .B(_4504__bF_buf1), .C(_4700_), .Y(_4701_) );
	NAND3X1 NAND3X1_994 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .B(_4701_), .C(_4699_), .Y(_4702_) );
	NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_4698_), .B(_4696_), .Y(_4703_) );
	NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_4703_), .B(divider_divuResult_11_bF_buf2), .Y(_4704_) );
	OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf4), .B(_4504__bF_buf0), .C(_4272_), .Y(_4705_) );
	NAND3X1 NAND3X1_995 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf1), .B(_4705_), .C(_4704_), .Y(_4706_) );
	AOI22X1 AOI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_4702_), .B(_4706_), .C(_4695_), .D(_4688_), .Y(_4707_) );
	NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_4707_), .B(_4677_), .Y(_4708_) );
	NAND3X1 NAND3X1_996 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(_4296_), .C(_4482_), .Y(_4709_) );
	NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_4291_), .B(_4297_), .Y(_4710_) );
	INVX1 INVX1_808 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .Y(_4711_) );
	OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_4711_), .B(_4409_), .C(_4452_), .Y(_4712_) );
	OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_4447_), .B(_4448_), .C(_4712_), .Y(_4713_) );
	NAND3X1 NAND3X1_997 ( .gnd(gnd), .vdd(vdd), .A(_4710_), .B(_4336_), .C(_4713_), .Y(_4715_) );
	NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_4303_), .B(_4307_), .Y(_4716_) );
	INVX1 INVX1_809 ( .gnd(gnd), .vdd(vdd), .A(_4716_), .Y(_4717_) );
	AOI21X1 AOI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_4418_), .C(_4329_), .Y(_4718_) );
	OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_4717_), .B(_4718_), .C(_4336_), .Y(_4719_) );
	OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_4330_), .B(_4334_), .C(_4719_), .Y(_4720_) );
	NAND3X1 NAND3X1_998 ( .gnd(gnd), .vdd(vdd), .A(_4715_), .B(_4720_), .C(divider_divuResult_11_bF_buf1), .Y(_4721_) );
	NAND3X1 NAND3X1_999 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_4709_), .C(_4721_), .Y(_4722_) );
	NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(_4296_), .Y(_4723_) );
	OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(_4723_), .Y(_4724_) );
	INVX1 INVX1_810 ( .gnd(gnd), .vdd(vdd), .A(_4710_), .Y(_4726_) );
	NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_4719_), .Y(_4727_) );
	AOI21X1 AOI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_4713_), .B(_4336_), .C(_4710_), .Y(_4728_) );
	OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_4728_), .B(_4727_), .C(divider_divuResult_11_bF_buf0), .Y(_4729_) );
	NAND3X1 NAND3X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf6), .B(_4724_), .C(_4729_), .Y(_4730_) );
	NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4278_), .Y(_4731_) );
	AOI21X1 AOI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_4731_), .C(_4350_), .Y(_4732_) );
	OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_4426_), .B(_4732_), .C(_4185_), .Y(_4733_) );
	NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_4717_), .B(_4718_), .Y(_4734_) );
	NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_4713_), .B(_4734_), .Y(_4735_) );
	NAND3X1 NAND3X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4735_), .C(_4733_), .Y(_4737_) );
	INVX1 INVX1_811 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .Y(_4738_) );
	OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf2), .B(_4504__bF_buf3), .C(_4738_), .Y(_4739_) );
	NAND3X1 NAND3X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf1), .B(_4739_), .C(_4737_), .Y(_4740_) );
	OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf1), .B(_4504__bF_buf2), .C(_4335_), .Y(_4741_) );
	AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_4734_), .B(_4713_), .Y(_4742_) );
	NAND3X1 NAND3X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4733_), .C(_4742_), .Y(_4743_) );
	NAND3X1 NAND3X1_1004 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_4741_), .C(_4743_), .Y(_4744_) );
	NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(_4744_), .Y(_4745_) );
	AOI21X1 AOI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .B(_4730_), .C(_4745_), .Y(_4746_) );
	OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf0), .B(_4504__bF_buf1), .C(_4321_), .Y(_4748_) );
	NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_4412_), .B(_4413_), .Y(_4749_) );
	AOI21X1 AOI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_4416_), .B(_4417_), .C(_4409_), .Y(_4750_) );
	OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .B(_4750_), .C(_4749_), .Y(_4751_) );
	INVX1 INVX1_812 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .Y(_4752_) );
	INVX1 INVX1_813 ( .gnd(gnd), .vdd(vdd), .A(_4749_), .Y(_4753_) );
	NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_4417_), .B(_4416_), .Y(_4754_) );
	NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_4754_), .B(_4479_), .Y(_4755_) );
	NAND3X1 NAND3X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_4752_), .B(_4753_), .C(_4755_), .Y(_4756_) );
	NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_4751_), .Y(_4757_) );
	OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4757_), .C(_4748_), .Y(_4759_) );
	NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf0), .B(_4759_), .Y(_4760_) );
	INVX1 INVX1_814 ( .gnd(gnd), .vdd(vdd), .A(_4321_), .Y(_4761_) );
	OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf4), .B(_4504__bF_buf0), .C(_4761_), .Y(_4762_) );
	NAND3X1 NAND3X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4757_), .C(_4733_), .Y(_4763_) );
	AOI21X1 AOI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .B(_4762_), .C(_4714__bF_buf6), .Y(_4764_) );
	NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_4754_), .B(_4479_), .Y(_4765_) );
	NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_4750_), .B(_4765_), .Y(_4766_) );
	INVX1 INVX1_815 ( .gnd(gnd), .vdd(vdd), .A(_4766_), .Y(_4767_) );
	NAND3X1 NAND3X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4767_), .C(_4733_), .Y(_4768_) );
	OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .B(divider_divuResult_12_bF_buf6), .C(_4325_), .Y(_4770_) );
	INVX1 INVX1_816 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .Y(_4771_) );
	OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(_4771_), .Y(_4772_) );
	NAND3X1 NAND3X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_4772_), .C(_4768_), .Y(_4773_) );
	OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_4773_), .B(_4764_), .C(_4760_), .Y(_4774_) );
	NAND3X1 NAND3X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf5), .B(_4709_), .C(_4721_), .Y(_4775_) );
	AOI21X1 AOI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_4721_), .B(_4709_), .C(_8971__bF_buf4), .Y(_4776_) );
	OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(_4776_), .C(_4775_), .Y(_4777_) );
	AOI21X1 AOI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_4746_), .B(_4774_), .C(_4777_), .Y(_4778_) );
	NAND3X1 NAND3X1_1010 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .B(_4665_), .C(_4664_), .Y(_4779_) );
	NAND3X1 NAND3X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf4), .B(_4687_), .C(_4678_), .Y(_4781_) );
	AOI21X1 AOI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_4678_), .B(_4687_), .C(_1265__bF_buf3), .Y(_4782_) );
	OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_4700_), .B(divider_divuResult_11_bF_buf5), .C(_4704_), .Y(_4783_) );
	NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf0), .B(_4783_), .Y(_4784_) );
	AOI21X1 AOI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_4784_), .B(_4781_), .C(_4782_), .Y(_4785_) );
	NAND3X1 NAND3X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf3), .B(_4645_), .C(_4659_), .Y(_4786_) );
	OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .B(divider_divuResult_11_bF_buf4), .C(_4668_), .Y(_4787_) );
	OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .B(_4787_), .C(_4786_), .Y(_4788_) );
	AOI22X1 AOI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_4779_), .B(_4788_), .C(_4785_), .D(_4677_), .Y(_4789_) );
	OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_4708_), .B(_4778_), .C(_4789_), .Y(_4790_) );
	NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_4476_), .B(_4469_), .Y(_4792_) );
	AOI21X1 AOI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf1), .B(_4405_), .C(_4474_), .Y(_4793_) );
	XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(_4792_), .Y(_4794_) );
	NAND3X1 NAND3X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4794_), .C(_4733_), .Y(_4795_) );
	OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf2), .B(_4504__bF_buf3), .C(_4389_), .Y(_4796_) );
	NAND3X1 NAND3X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_4796_), .C(_4795_), .Y(_4797_) );
	INVX1 INVX1_817 ( .gnd(gnd), .vdd(vdd), .A(_4794_), .Y(_4798_) );
	NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf1), .B(_4798_), .C(_4504__bF_buf2), .Y(_4799_) );
	AOI22X1 AOI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_4388_), .C(_4009_), .D(_4733_), .Y(_4800_) );
	OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_4799_), .B(_4800_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .Y(_4801_) );
	NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(_4801_), .Y(_4803_) );
	NAND3X1 NAND3X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .B(_4471_), .C(_4472_), .Y(_4804_) );
	AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_4804_), .B(_4403_), .Y(_4805_) );
	INVX1 INVX1_818 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .Y(_4806_) );
	NAND3X1 NAND3X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4806_), .C(_4733_), .Y(_4807_) );
	OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf0), .B(_4504__bF_buf1), .C(_4475_), .Y(_4808_) );
	NAND3X1 NAND3X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_4808_), .C(_4807_), .Y(_4809_) );
	OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf4), .B(_4504__bF_buf0), .C(_4405_), .Y(_4810_) );
	NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .B(divider_divuResult_11_bF_buf3), .Y(_4811_) );
	NAND3X1 NAND3X1_1018 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .B(_4810_), .C(_4811_), .Y(_4812_) );
	NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(_4812_), .Y(_4814_) );
	NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(_4470_), .Y(_4815_) );
	NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .B(_4815_), .Y(_4816_) );
	INVX1 INVX1_819 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .Y(_4817_) );
	NAND3X1 NAND3X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4817_), .C(_4733_), .Y(_4818_) );
	OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(divider_aOp_abs_11_), .Y(_4819_) );
	AOI21X1 AOI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .B(_4819_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .Y(_4820_) );
	NAND3X1 NAND3X1_1020 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .B(_4819_), .C(_4818_), .Y(_4821_) );
	NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_10_), .B(_1746__bF_buf1), .Y(_4822_) );
	INVX1 INVX1_820 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .Y(_4823_) );
	AOI21X1 AOI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_4821_), .B(_4823_), .C(_4820_), .Y(_4825_) );
	NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4814_), .B(_4803_), .C(_4825_), .Y(_4826_) );
	OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_4059_), .B(divider_divuResult_12_bF_buf5), .C(_4359_), .Y(_4827_) );
	OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf2), .B(_4504__bF_buf3), .C(_4827_), .Y(_4828_) );
	INVX1 INVX1_821 ( .gnd(gnd), .vdd(vdd), .A(_4467_), .Y(_4829_) );
	OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_4829_), .B(_4478_), .C(_4369_), .Y(_4830_) );
	XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_4830_), .B(_4374_), .Y(_4831_) );
	NAND3X1 NAND3X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4831_), .C(_4733_), .Y(_4832_) );
	NAND3X1 NAND3X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf1), .B(_4828_), .C(_4832_), .Y(_4833_) );
	INVX1 INVX1_822 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .Y(_4834_) );
	NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_4467_), .B(_4407_), .Y(_4836_) );
	NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_4829_), .B(_4478_), .Y(_4837_) );
	NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_4836_), .B(_4837_), .Y(_4838_) );
	INVX1 INVX1_823 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .Y(_4839_) );
	NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_4839_), .B(divider_divuResult_11_bF_buf2), .Y(_4840_) );
	OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf1), .B(_4504__bF_buf2), .C(_4368_), .Y(_4841_) );
	AOI21X1 AOI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(_4841_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .Y(_4842_) );
	INVX1 INVX1_824 ( .gnd(gnd), .vdd(vdd), .A(_4831_), .Y(_4843_) );
	OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4843_), .C(_4828_), .Y(_4844_) );
	NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .B(_4844_), .Y(_4845_) );
	AOI21X1 AOI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_4845_), .B(_4842_), .C(_4834_), .Y(_4847_) );
	NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_4799_), .B(_4800_), .Y(_4848_) );
	OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4805_), .C(_4808_), .Y(_4849_) );
	OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_4849_), .C(_4797_), .Y(_4850_) );
	OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_4848_), .C(_4850_), .Y(_4851_) );
	NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(_4851_), .Y(_4852_) );
	NAND3X1 NAND3X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4838_), .C(_4733_), .Y(_4853_) );
	OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf0), .B(_4504__bF_buf1), .C(_4464_), .Y(_4854_) );
	NAND3X1 NAND3X1_1024 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .B(_4854_), .C(_4853_), .Y(_4855_) );
	NAND3X1 NAND3X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_4841_), .C(_4840_), .Y(_4856_) );
	NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_4855_), .B(_4856_), .Y(_4858_) );
	NAND3X1 NAND3X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_4833_), .B(_4845_), .C(_4858_), .Y(_4859_) );
	NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(_4859_), .Y(_4860_) );
	OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_4852_), .B(_4826_), .C(_4860_), .Y(_4861_) );
	NAND3X1 NAND3X1_1027 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .B(_4724_), .C(_4729_), .Y(_4862_) );
	NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_4775_), .B(_4862_), .Y(_4863_) );
	NAND3X1 NAND3X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_4752_), .B(_4749_), .C(_4755_), .Y(_4864_) );
	OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .B(_4750_), .C(_4753_), .Y(_4865_) );
	NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .B(_4865_), .Y(_4866_) );
	NAND3X1 NAND3X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4866_), .C(_4733_), .Y(_4867_) );
	AOI21X1 AOI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_4867_), .B(_4748_), .C(_4714__bF_buf5), .Y(_4869_) );
	AOI21X1 AOI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .B(_4762_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .Y(_4870_) );
	NAND3X1 NAND3X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4766_), .C(_4733_), .Y(_4871_) );
	OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf4), .B(_4504__bF_buf0), .C(_4770_), .Y(_4872_) );
	AOI21X1 AOI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_4871_), .B(_4872_), .C(_4999__bF_buf3), .Y(_4873_) );
	AOI21X1 AOI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_4768_), .B(_4772_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .Y(_4874_) );
	OAI22X1 OAI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_4873_), .B(_4874_), .C(_4869_), .D(_4870_), .Y(_4875_) );
	NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(_4863_), .C(_4875_), .Y(_4876_) );
	NAND3X1 NAND3X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_4677_), .B(_4707_), .C(_4876_), .Y(_4877_) );
	NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_4877_), .B(_4861_), .Y(_4878_) );
	OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_4878_), .C(_4644_), .Y(_4880_) );
	AOI21X1 AOI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .B(_4615_), .C(_2097_), .Y(divider_divuResult_10_) );
	INVX8 INVX8_36 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf1), .Y(_4881_) );
	INVX1 INVX1_825 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .Y(_4882_) );
	INVX1 INVX1_826 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .Y(_4883_) );
	AOI22X1 AOI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_4573_), .C(_4883_), .D(_4882_), .Y(_4884_) );
	NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_4486_), .Y(_4885_) );
	AOI21X1 AOI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_4618_), .C(_4885_), .Y(_4886_) );
	INVX1 INVX1_827 ( .gnd(gnd), .vdd(vdd), .A(_4533_), .Y(_4887_) );
	AOI21X1 AOI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_4527_), .B(_4538_), .C(_4887_), .Y(_4888_) );
	OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_4885_), .B(_4507_), .C(_4486_), .Y(_4890_) );
	AOI21X1 AOI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4886_), .C(_4890_), .Y(_4891_) );
	OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_4624_), .B(_4884_), .C(_4891_), .Y(_4892_) );
	NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_4642_), .B(_4585_), .Y(_4893_) );
	NAND3X1 NAND3X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_4623_), .B(_4886_), .C(_4893_), .Y(_4894_) );
	NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_4670_), .Y(_4895_) );
	NAND3X1 NAND3X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_4786_), .B(_4779_), .C(_4895_), .Y(_4896_) );
	NAND3X1 NAND3X1_1034 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .B(_4689_), .C(_4694_), .Y(_4897_) );
	NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_4706_), .B(_4702_), .Y(_4898_) );
	NAND3X1 NAND3X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_4781_), .B(_4897_), .C(_4898_), .Y(_4899_) );
	NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .B(_4896_), .Y(_4901_) );
	NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .B(_4730_), .Y(_4902_) );
	AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_4744_), .B(_4740_), .Y(_4903_) );
	NAND3X1 NAND3X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .B(_4902_), .C(_4774_), .Y(_4904_) );
	INVX1 INVX1_828 ( .gnd(gnd), .vdd(vdd), .A(_4775_), .Y(_4905_) );
	INVX1 INVX1_829 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .Y(_4906_) );
	AOI21X1 AOI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_4906_), .B(_4862_), .C(_4905_), .Y(_4907_) );
	NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_4907_), .B(_4904_), .Y(_4908_) );
	AOI21X1 AOI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .B(_4689_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .Y(_4909_) );
	AOI21X1 AOI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4705_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .Y(_4910_) );
	OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .B(_4909_), .C(_4897_), .Y(_4912_) );
	AOI21X1 AOI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_4664_), .B(_4665_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .Y(_4913_) );
	AOI21X1 AOI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_4675_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .Y(_4914_) );
	OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_4914_), .B(_4913_), .C(_4779_), .Y(_4915_) );
	OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_4912_), .B(_4896_), .C(_4915_), .Y(_4916_) );
	AOI21X1 AOI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(_4908_), .C(_4916_), .Y(_4917_) );
	AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(_4797_), .Y(_4918_) );
	NAND3X1 NAND3X1_1037 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_4808_), .C(_4807_), .Y(_4919_) );
	NAND3X1 NAND3X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_4810_), .C(_4811_), .Y(_4920_) );
	NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(_4920_), .Y(_4921_) );
	NAND3X1 NAND3X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4816_), .C(_4733_), .Y(_4923_) );
	OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_4010__bF_buf3), .B(_4504__bF_buf4), .C(_4470_), .Y(_4924_) );
	NAND3X1 NAND3X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf0), .B(_4924_), .C(_4923_), .Y(_4925_) );
	AOI21X1 AOI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_4923_), .B(_4924_), .C(_1768__bF_buf7), .Y(_4926_) );
	OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .B(_4926_), .C(_4925_), .Y(_4927_) );
	NAND3X1 NAND3X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_4921_), .B(_4927_), .C(_4918_), .Y(_4928_) );
	NAND3X1 NAND3X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf7), .B(_4854_), .C(_4853_), .Y(_4929_) );
	AOI21X1 AOI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_4828_), .C(_4100__bF_buf0), .Y(_4930_) );
	OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_4929_), .B(_4930_), .C(_4833_), .Y(_4931_) );
	AOI21X1 AOI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_4850_), .B(_4801_), .C(_4931_), .Y(_4932_) );
	AOI22X1 AOI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(_4859_), .C(_4932_), .D(_4928_), .Y(_4934_) );
	NAND3X1 NAND3X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(_4876_), .C(_4934_), .Y(_4935_) );
	AOI21X1 AOI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_4917_), .C(_4894_), .Y(_4936_) );
	OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_4936_), .C(_3171__bF_buf2), .Y(_4937_) );
	AOI21X1 AOI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_4937__bF_buf5), .B(_4485_), .C(_2240__bF_buf4), .Y(_4938_) );
	XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(_4881__bF_buf3), .Y(_4939_) );
	INVX1 INVX1_830 ( .gnd(gnd), .vdd(vdd), .A(_4619_), .Y(_4940_) );
	AOI21X1 AOI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_4917_), .C(_4643_), .Y(_4941_) );
	OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_4607_), .B(_4941_), .C(_4623_), .Y(_4942_) );
	AOI21X1 AOI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_4942_), .B(_4610_), .C(_4940_), .Y(_4943_) );
	NAND3X1 NAND3X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_4940_), .B(_4610_), .C(_4942_), .Y(_4945_) );
	INVX1 INVX1_831 ( .gnd(gnd), .vdd(vdd), .A(_4945_), .Y(_4946_) );
	OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4946_), .C(divider_divuResult_10_bF_buf5), .Y(_4947_) );
	OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_4503_), .B(divider_divuResult_11_bF_buf1), .C(_4510_), .Y(_4948_) );
	OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf4), .B(_4948_), .Y(_4949_) );
	NAND3X1 NAND3X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf2), .B(_4949_), .C(_4947_), .Y(_4950_) );
	NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_4610_), .B(_4942_), .Y(_4951_) );
	NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_4619_), .B(_4951_), .Y(_4952_) );
	NAND3X1 NAND3X1_1046 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf3), .B(_4945_), .C(_4952_), .Y(_4953_) );
	NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_4948_), .B(_4937__bF_buf4), .Y(_4954_) );
	NAND3X1 NAND3X1_1047 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf3), .B(_4954_), .C(_4953_), .Y(_4956_) );
	NAND3X1 NAND3X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_4939_), .B(_4956_), .C(_4950_), .Y(_4957_) );
	OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(divider_divuResult_11_bF_buf0), .C(_4531_), .Y(_4958_) );
	NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_4958_), .B(divider_divuResult_10_bF_buf2), .Y(_4959_) );
	INVX1 INVX1_832 ( .gnd(gnd), .vdd(vdd), .A(_4959_), .Y(_4960_) );
	NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4621_), .Y(_4961_) );
	INVX1 INVX1_833 ( .gnd(gnd), .vdd(vdd), .A(_4961_), .Y(_4962_) );
	OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_4607_), .B(_4941_), .C(_4543_), .Y(_4963_) );
	AOI21X1 AOI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4538_), .C(_4962_), .Y(_4964_) );
	NAND3X1 NAND3X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_4962_), .B(_4538_), .C(_4963_), .Y(_4965_) );
	INVX1 INVX1_834 ( .gnd(gnd), .vdd(vdd), .A(_4965_), .Y(_4967_) );
	OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_4964_), .B(_4967_), .C(divider_divuResult_10_bF_buf1), .Y(_4968_) );
	NAND3X1 NAND3X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf0), .B(_4960_), .C(_4968_), .Y(_4969_) );
	OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_4878_), .C(_4893_), .Y(_4970_) );
	AOI21X1 AOI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_4970_), .B(_4884_), .C(_4622_), .Y(_4971_) );
	OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_4609_), .B(_4971_), .C(_4961_), .Y(_4972_) );
	AOI21X1 AOI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_4972_), .B(_4965_), .C(_4937__bF_buf3), .Y(_4973_) );
	OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_4959_), .B(_4973_), .C(divider_absoluteValue_B_flipSign_result_20_bF_buf0), .Y(_4974_) );
	NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_4543_), .B(_4607_), .C(_4941_), .Y(_4975_) );
	OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_4975_), .B(_4971_), .C(divider_divuResult_10_bF_buf0), .Y(_4976_) );
	OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_4180_), .B(divider_divuResult_11_bF_buf5), .C(_4536_), .Y(_4978_) );
	NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_4978_), .B(_4937__bF_buf2), .Y(_4979_) );
	NAND3X1 NAND3X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf4), .B(_4979_), .C(_4976_), .Y(_4980_) );
	NAND3X1 NAND3X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_4536_), .B(_4537_), .C(_4937__bF_buf1), .Y(_4981_) );
	NAND3X1 NAND3X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_4622_), .B(_4884_), .C(_4970_), .Y(_4982_) );
	NAND3X1 NAND3X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4982_), .C(divider_divuResult_10_bF_buf5), .Y(_4983_) );
	NAND3X1 NAND3X1_1055 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf4), .B(_4981_), .C(_4983_), .Y(_4984_) );
	AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_4980_), .B(_4984_), .Y(_4985_) );
	NAND3X1 NAND3X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_4985_), .B(_4969_), .C(_4974_), .Y(_4986_) );
	NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_4957_), .B(_4986_), .Y(_4987_) );
	NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_4937__bF_buf0), .Y(_4989_) );
	NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf2), .B(_4571_), .Y(_4990_) );
	NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_4567_), .Y(_4991_) );
	INVX1 INVX1_835 ( .gnd(gnd), .vdd(vdd), .A(_4991_), .Y(_4992_) );
	INVX1 INVX1_836 ( .gnd(gnd), .vdd(vdd), .A(_4584_), .Y(_4993_) );
	INVX1 INVX1_837 ( .gnd(gnd), .vdd(vdd), .A(_4642_), .Y(_4994_) );
	OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .B(_4878_), .C(_4994_), .Y(_4995_) );
	AOI21X1 AOI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_4995_), .B(_4606_), .C(_4993_), .Y(_4996_) );
	OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_4990_), .B(_4996_), .C(_4992_), .Y(_4997_) );
	INVX1 INVX1_838 ( .gnd(gnd), .vdd(vdd), .A(_4990_), .Y(_4998_) );
	AOI21X1 AOI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_4917_), .C(_4642_), .Y(_5000_) );
	OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_4883_), .B(_5000_), .C(_4584_), .Y(_5001_) );
	NAND3X1 NAND3X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(_4991_), .C(_5001_), .Y(_5002_) );
	NAND3X1 NAND3X1_1058 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf4), .B(_5002_), .C(_4997_), .Y(_5003_) );
	NAND3X1 NAND3X1_1059 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf1), .B(_4989_), .C(_5003_), .Y(_5004_) );
	INVX1 INVX1_839 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .Y(_5005_) );
	OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf3), .B(_4562_), .Y(_5006_) );
	NAND3X1 NAND3X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(_4992_), .C(_5001_), .Y(_5007_) );
	OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_4990_), .B(_4996_), .C(_4991_), .Y(_5008_) );
	NAND3X1 NAND3X1_1061 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf2), .B(_5007_), .C(_5008_), .Y(_5009_) );
	NAND3X1 NAND3X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf1), .B(_5006_), .C(_5009_), .Y(_5011_) );
	INVX1 INVX1_840 ( .gnd(gnd), .vdd(vdd), .A(_4571_), .Y(_5012_) );
	NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_5012_), .B(_4937__bF_buf5), .Y(_5013_) );
	NAND3X1 NAND3X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_4993_), .B(_4606_), .C(_4995_), .Y(_5014_) );
	NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_5014_), .Y(_5015_) );
	OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_4937__bF_buf4), .B(_5015_), .C(_5013_), .Y(_5016_) );
	NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf3), .B(_5016_), .Y(_5017_) );
	AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_5011_), .B(_5017_), .Y(_5018_) );
	NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .B(_5016_), .Y(_5019_) );
	NAND3X1 NAND3X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_5014_), .C(divider_divuResult_10_bF_buf1), .Y(_5020_) );
	NAND3X1 NAND3X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf2), .B(_5013_), .C(_5020_), .Y(_5022_) );
	NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_5022_), .B(_5019_), .Y(_5023_) );
	NAND3X1 NAND3X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(_5011_), .C(_5023_), .Y(_5024_) );
	INVX1 INVX1_841 ( .gnd(gnd), .vdd(vdd), .A(_4603_), .Y(_5025_) );
	NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_4634_), .Y(_5026_) );
	INVX1 INVX1_842 ( .gnd(gnd), .vdd(vdd), .A(_4641_), .Y(_5027_) );
	INVX1 INVX1_843 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .Y(_5028_) );
	NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_4746_), .B(_5028_), .Y(_5029_) );
	NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(_4708_), .Y(_5030_) );
	AOI21X1 AOI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_5030_), .C(_4790_), .Y(_5031_) );
	NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_5027_), .B(_5031_), .Y(_5033_) );
	OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .B(_5033_), .C(_5026_), .Y(_5034_) );
	INVX1 INVX1_844 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .Y(_5035_) );
	NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .B(_5033_), .Y(_5036_) );
	NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_5035_), .B(_5036_), .Y(_5037_) );
	NAND3X1 NAND3X1_1067 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf0), .B(_5034_), .C(_5037_), .Y(_5038_) );
	NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_4599_), .B(_4937__bF_buf3), .Y(_5039_) );
	NAND3X1 NAND3X1_1068 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf1), .B(_5039_), .C(_5038_), .Y(_5040_) );
	AOI21X1 AOI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_5038_), .B(_5039_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf0), .Y(_5041_) );
	AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_5031_), .B(_5027_), .Y(_5042_) );
	OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_5033_), .B(_5042_), .C(divider_divuResult_10_bF_buf5), .Y(_5044_) );
	NAND3X1 NAND3X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_4639_), .C(_4937__bF_buf2), .Y(_5045_) );
	NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_5045_), .B(_5044_), .Y(_5046_) );
	NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .B(_5046_), .Y(_5047_) );
	OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(_5041_), .C(_5040_), .Y(_5048_) );
	OAI22X1 OAI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_5005_), .B(_5018_), .C(_5048_), .D(_5024_), .Y(_5049_) );
	NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf3), .B(_4959_), .C(_4973_), .Y(_5050_) );
	INVX1 INVX1_845 ( .gnd(gnd), .vdd(vdd), .A(_4980_), .Y(_5051_) );
	AOI21X1 AOI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_4974_), .B(_5051_), .C(_5050_), .Y(_5052_) );
	NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf0), .B(_4938_), .Y(_5053_) );
	AOI21X1 AOI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_4953_), .B(_4954_), .C(divider_absoluteValue_B_flipSign_result_21_bF_buf2), .Y(_5055_) );
	AOI21X1 AOI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_5055_), .B(_4939_), .C(_5053_), .Y(_5056_) );
	OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_4957_), .B(_5052_), .C(_5056_), .Y(_5057_) );
	AOI21X1 AOI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_5049_), .C(_5057_), .Y(_5058_) );
	AOI21X1 AOI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_5038_), .B(_5039_), .C(_2922__bF_buf2), .Y(_5059_) );
	NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_4598_), .B(_4937__bF_buf1), .Y(_5060_) );
	OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .B(_5033_), .C(_5035_), .Y(_5061_) );
	OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_4629_), .B(_4635_), .C(_5036_), .Y(_5062_) );
	NAND3X1 NAND3X1_1070 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf4), .B(_5061_), .C(_5062_), .Y(_5063_) );
	AOI21X1 AOI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_5063_), .B(_5060_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .Y(_5064_) );
	NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf3), .B(_5046_), .Y(_5066_) );
	AOI21X1 AOI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_5044_), .B(_5045_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .Y(_5067_) );
	OAI22X1 OAI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_5066_), .B(_5067_), .C(_5059_), .D(_5064_), .Y(_5068_) );
	NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_5068_), .B(_5024_), .Y(_5069_) );
	OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_4458_), .B(divider_divuResult_11_bF_buf4), .C(_4659_), .Y(_5070_) );
	INVX1 INVX1_846 ( .gnd(gnd), .vdd(vdd), .A(_5070_), .Y(_5071_) );
	NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_5071_), .B(_4937__bF_buf0), .Y(_5072_) );
	NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_4661_), .B(_4666_), .Y(_5073_) );
	INVX1 INVX1_847 ( .gnd(gnd), .vdd(vdd), .A(_4914_), .Y(_5074_) );
	INVX1 INVX1_848 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .Y(_5075_) );
	OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(divider_divuResult_11_bF_buf3), .C(_4687_), .Y(_5077_) );
	OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .B(_5077_), .C(_4784_), .Y(_5078_) );
	OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(_4861_), .C(_4778_), .Y(_5079_) );
	AOI22X1 AOI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .B(_5078_), .C(_4707_), .D(_5079_), .Y(_5080_) );
	OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .B(_5080_), .C(_5074_), .Y(_5081_) );
	NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .B(_5081_), .Y(_5082_) );
	INVX1 INVX1_849 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .Y(_5083_) );
	AOI21X1 AOI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_4876_), .C(_4908_), .Y(_5084_) );
	OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .B(_5084_), .C(_4912_), .Y(_5085_) );
	NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .B(_5085_), .Y(_5086_) );
	NAND3X1 NAND3X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_5074_), .C(_5086_), .Y(_5088_) );
	NAND3X1 NAND3X1_1072 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf3), .B(_5088_), .C(_5082_), .Y(_5089_) );
	NAND3X1 NAND3X1_1073 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf0), .B(_5072_), .C(_5089_), .Y(_5090_) );
	AOI21X1 AOI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .B(_5072_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .Y(_5091_) );
	NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .B(_5080_), .Y(_5092_) );
	NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .B(_5085_), .Y(_5093_) );
	OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .B(_5092_), .C(divider_divuResult_10_bF_buf2), .Y(_5094_) );
	NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_4787_), .B(_4937__bF_buf5), .Y(_5095_) );
	NAND3X1 NAND3X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf2), .B(_5095_), .C(_5094_), .Y(_5096_) );
	INVX1 INVX1_850 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .Y(_5097_) );
	OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .B(_5091_), .C(_5090_), .Y(_5099_) );
	NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_5070_), .B(_4937__bF_buf4), .Y(_5100_) );
	NAND3X1 NAND3X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .B(_5074_), .C(_5086_), .Y(_5101_) );
	NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_5081_), .Y(_5102_) );
	NAND3X1 NAND3X1_1076 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf1), .B(_5101_), .C(_5102_), .Y(_5103_) );
	NAND3X1 NAND3X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf0), .B(_5100_), .C(_5103_), .Y(_5104_) );
	NAND3X1 NAND3X1_1078 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .B(_5095_), .C(_5094_), .Y(_5105_) );
	NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .B(_5080_), .Y(_5106_) );
	AOI21X1 AOI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5086_), .C(_4937__bF_buf3), .Y(_5107_) );
	AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_4937__bF_buf2), .B(_4787_), .Y(_5108_) );
	OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .B(_5107_), .C(_1494__bF_buf1), .Y(_5110_) );
	NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_5110_), .Y(_5111_) );
	NAND3X1 NAND3X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .B(_5090_), .C(_5111_), .Y(_5112_) );
	INVX1 INVX1_851 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .Y(_5113_) );
	NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(divider_divuResult_10_bF_buf0), .Y(_5114_) );
	NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_4695_), .B(_4688_), .Y(_5115_) );
	INVX1 INVX1_852 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .Y(_5116_) );
	OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_5084_), .C(_4784_), .Y(_5117_) );
	NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .B(_5117_), .Y(_5118_) );
	INVX1 INVX1_853 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .Y(_5119_) );
	NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_5079_), .Y(_5121_) );
	NAND3X1 NAND3X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_4784_), .C(_5121_), .Y(_5122_) );
	AOI21X1 AOI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .B(_5118_), .C(_4937__bF_buf1), .Y(_5123_) );
	OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .B(_5114_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .Y(_5124_) );
	NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .B(_5123_), .C(_5114_), .Y(_5125_) );
	OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_4894_), .B(_5031_), .C(_4615_), .Y(_5126_) );
	NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_5084_), .Y(_5127_) );
	NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .B(_5121_), .Y(_5128_) );
	NAND3X1 NAND3X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf1), .B(_5126__bF_buf3), .C(_5128_), .Y(_5129_) );
	NAND3X1 NAND3X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4705_), .C(_4937__bF_buf0), .Y(_5130_) );
	NAND3X1 NAND3X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf2), .B(_5129_), .C(_5130_), .Y(_5132_) );
	INVX1 INVX1_854 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .Y(_5133_) );
	OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_5125_), .C(_5124_), .Y(_5134_) );
	OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_5134_), .B(_5112_), .C(_5099_), .Y(_5135_) );
	NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .B(divider_divuResult_10_bF_buf5), .Y(_5136_) );
	NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .B(_5122_), .Y(_5137_) );
	NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_4937__bF_buf5), .B(_5137_), .Y(_5138_) );
	OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5138_), .C(_1484__bF_buf1), .Y(_5139_) );
	NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(_4937__bF_buf4), .Y(_5140_) );
	XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .B(_4898_), .Y(_5141_) );
	NAND3X1 NAND3X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf0), .B(_5126__bF_buf2), .C(_5141_), .Y(_5143_) );
	NAND3X1 NAND3X1_1085 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .B(_5143_), .C(_5140_), .Y(_5144_) );
	AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_5144_), .Y(_5145_) );
	NAND3X1 NAND3X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_5124_), .B(_5139_), .C(_5145_), .Y(_5146_) );
	NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_5146_), .B(_5112_), .Y(_5147_) );
	NAND3X1 NAND3X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_4724_), .B(_4729_), .C(_4937__bF_buf3), .Y(_5148_) );
	AOI21X1 AOI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_5028_), .C(_4774_), .Y(_5149_) );
	OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(_5149_), .C(_4740_), .Y(_5150_) );
	AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_5150_), .B(_4902_), .Y(_5151_) );
	NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_4902_), .B(_5150_), .Y(_5152_) );
	OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_5152_), .B(_5151_), .C(divider_divuResult_10_bF_buf4), .Y(_5154_) );
	NAND3X1 NAND3X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf5), .B(_5148_), .C(_5154_), .Y(_5155_) );
	INVX1 INVX1_855 ( .gnd(gnd), .vdd(vdd), .A(_5155_), .Y(_5156_) );
	NAND3X1 NAND3X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(_4721_), .C(_4937__bF_buf2), .Y(_5157_) );
	NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_4902_), .B(_5150_), .Y(_5158_) );
	OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_5150_), .B(_4902_), .Y(_5159_) );
	NAND3X1 NAND3X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_5159_), .C(divider_divuResult_10_bF_buf3), .Y(_5160_) );
	NAND3X1 NAND3X1_1091 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .B(_5157_), .C(_5160_), .Y(_5161_) );
	XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_5149_), .B(_4903_), .Y(_5162_) );
	NAND3X1 NAND3X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf3), .B(_5126__bF_buf1), .C(_5162_), .Y(_5163_) );
	OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4735_), .C(_4741_), .Y(_5165_) );
	NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_5165_), .B(_4937__bF_buf1), .Y(_5166_) );
	AOI21X1 AOI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_5166_), .B(_5163_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .Y(_5167_) );
	AOI21X1 AOI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_5161_), .B(_5167_), .C(_5156_), .Y(_5168_) );
	XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_5149_), .B(_4745_), .Y(_5169_) );
	NAND3X1 NAND3X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf2), .B(_5126__bF_buf0), .C(_5169_), .Y(_5170_) );
	INVX1 INVX1_856 ( .gnd(gnd), .vdd(vdd), .A(_5165_), .Y(_5171_) );
	NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_5171_), .B(_4937__bF_buf0), .Y(_5172_) );
	NAND3X1 NAND3X1_1094 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .B(_5170_), .C(_5172_), .Y(_5173_) );
	NAND3X1 NAND3X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf3), .B(_5163_), .C(_5166_), .Y(_5174_) );
	NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_5173_), .Y(_5176_) );
	NAND3X1 NAND3X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_5155_), .B(_5161_), .C(_5176_), .Y(_5177_) );
	NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_4759_), .Y(_5178_) );
	NAND3X1 NAND3X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf4), .B(_4748_), .C(_4867_), .Y(_5179_) );
	NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_5179_), .B(_5178_), .Y(_5180_) );
	INVX1 INVX1_857 ( .gnd(gnd), .vdd(vdd), .A(_4773_), .Y(_5181_) );
	INVX1 INVX1_858 ( .gnd(gnd), .vdd(vdd), .A(_4873_), .Y(_5182_) );
	INVX1 INVX1_859 ( .gnd(gnd), .vdd(vdd), .A(_4874_), .Y(_5183_) );
	NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_5182_), .B(_5183_), .Y(_5184_) );
	AOI21X1 AOI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_5184_), .C(_5181_), .Y(_5185_) );
	XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_5185_), .B(_5180_), .Y(_5187_) );
	NAND3X1 NAND3X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf1), .B(_5126__bF_buf3), .C(_5187_), .Y(_5188_) );
	OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_4759_), .B(divider_divuResult_10_bF_buf2), .C(_5188_), .Y(_5189_) );
	NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_5189_), .Y(_5190_) );
	NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .B(_5189_), .Y(_5191_) );
	OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4766_), .C(_4772_), .Y(_5192_) );
	INVX1 INVX1_860 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .Y(_5193_) );
	NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_5193_), .B(_4937__bF_buf5), .Y(_5194_) );
	XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_4934_), .B(_5184_), .Y(_5195_) );
	NAND3X1 NAND3X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf0), .B(_5195_), .C(_5126__bF_buf2), .Y(_5196_) );
	AOI21X1 AOI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_5194_), .B(_5196_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .Y(_5198_) );
	AOI21X1 AOI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(_5191_), .C(_5190_), .Y(_5199_) );
	OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_5199_), .B(_5177_), .C(_5168_), .Y(_5200_) );
	AOI21X1 AOI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_5147_), .B(_5200_), .C(_5135_), .Y(_5201_) );
	NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_4844_), .B(_4937__bF_buf4), .Y(_5202_) );
	NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_4930_), .B(_4834_), .Y(_5203_) );
	AOI22X1 AOI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_4855_), .B(_4856_), .C(_4851_), .D(_4928_), .Y(_5204_) );
	OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_4842_), .B(_5204_), .C(_5203_), .Y(_5205_) );
	NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_4842_), .B(_5204_), .Y(_5206_) );
	OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_4834_), .B(_4930_), .C(_5206_), .Y(_5207_) );
	NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_5205_), .B(_5207_), .Y(_5209_) );
	NAND3X1 NAND3X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf3), .B(_5209_), .C(_5126__bF_buf1), .Y(_5210_) );
	NAND3X1 NAND3X1_1101 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .B(_5210_), .C(_5202_), .Y(_5211_) );
	INVX1 INVX1_861 ( .gnd(gnd), .vdd(vdd), .A(_4844_), .Y(_5212_) );
	AOI21X1 AOI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_5126__bF_buf0), .B(_3171__bF_buf2), .C(_5212_), .Y(_5213_) );
	AOI21X1 AOI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_5205_), .B(_5207_), .C(_4937__bF_buf3), .Y(_5214_) );
	OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_5213_), .B(_5214_), .C(_4999__bF_buf2), .Y(_5215_) );
	NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(_4928_), .Y(_5216_) );
	NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(_5216_), .Y(_5217_) );
	NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_5204_), .B(_5217_), .Y(_5218_) );
	INVX1 INVX1_862 ( .gnd(gnd), .vdd(vdd), .A(_5218_), .Y(_5220_) );
	NAND3X1 NAND3X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf1), .B(_5220_), .C(_5126__bF_buf3), .Y(_5221_) );
	OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4839_), .C(_4854_), .Y(_5222_) );
	NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_5222_), .B(_4937__bF_buf2), .Y(_5223_) );
	NAND3X1 NAND3X1_1103 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_5221_), .C(_5223_), .Y(_5224_) );
	NAND3X1 NAND3X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf0), .B(_5218_), .C(_5126__bF_buf2), .Y(_5225_) );
	INVX1 INVX1_863 ( .gnd(gnd), .vdd(vdd), .A(_5222_), .Y(_5226_) );
	NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_5226_), .B(_4937__bF_buf1), .Y(_5227_) );
	NAND3X1 NAND3X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf7), .B(_5225_), .C(_5227_), .Y(_5228_) );
	AOI22X1 AOI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_5224_), .B(_5228_), .C(_5211_), .D(_5215_), .Y(_5229_) );
	OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_4814_), .B(_4825_), .C(_4809_), .Y(_5231_) );
	NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_4918_), .B(_5231_), .Y(_5232_) );
	OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_5231_), .B(_4918_), .Y(_5233_) );
	NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_5232_), .B(_5233_), .Y(_5234_) );
	NAND3X1 NAND3X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf3), .B(_5234_), .C(_5126__bF_buf1), .Y(_5235_) );
	INVX1 INVX1_864 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .Y(_5236_) );
	NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_5236_), .B(_4937__bF_buf0), .Y(_5237_) );
	NAND3X1 NAND3X1_1107 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .B(_5235_), .C(_5237_), .Y(_5238_) );
	AOI21X1 AOI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_5232_), .B(_5233_), .C(_4937__bF_buf5), .Y(_5239_) );
	AOI21X1 AOI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_5126__bF_buf0), .B(_3171__bF_buf2), .C(_4848_), .Y(_5240_) );
	OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_5240_), .B(_5239_), .C(_1735__bF_buf6), .Y(_5242_) );
	XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_4825_), .B(_4921_), .Y(_5243_) );
	INVX1 INVX1_865 ( .gnd(gnd), .vdd(vdd), .A(_5243_), .Y(_5244_) );
	NAND3X1 NAND3X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf1), .B(_5244_), .C(_5126__bF_buf3), .Y(_5245_) );
	NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_4849_), .B(_4937__bF_buf4), .Y(_5246_) );
	NAND3X1 NAND3X1_1109 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .B(_5245_), .C(_5246_), .Y(_5247_) );
	NAND3X1 NAND3X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf0), .B(_5243_), .C(_5126__bF_buf2), .Y(_5248_) );
	INVX1 INVX1_866 ( .gnd(gnd), .vdd(vdd), .A(_4849_), .Y(_5249_) );
	NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_5249_), .B(_4937__bF_buf3), .Y(_5250_) );
	NAND3X1 NAND3X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_5248_), .C(_5250_), .Y(_5251_) );
	AOI22X1 AOI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_5247_), .B(_5251_), .C(_5238_), .D(_5242_), .Y(_5253_) );
	NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_5229_), .B(_5253_), .Y(_5254_) );
	INVX1 INVX1_867 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_10_), .Y(_5255_) );
	NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(_5255_), .Y(_5256_) );
	NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .B(_5256_), .Y(_5257_) );
	NAND3X1 NAND3X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf3), .B(_5257_), .C(_5126__bF_buf1), .Y(_5258_) );
	NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_4937__bF_buf2), .Y(_5259_) );
	NAND3X1 NAND3X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf6), .B(_5258_), .C(_5259_), .Y(_5260_) );
	INVX1 INVX1_868 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .Y(_5261_) );
	NAND3X1 NAND3X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf2), .B(_5261_), .C(_5126__bF_buf0), .Y(_5262_) );
	NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_10_), .B(_4937__bF_buf1), .Y(_5264_) );
	NAND3X1 NAND3X1_1115 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_5262_), .C(_5264_), .Y(_5265_) );
	AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_5260_), .B(_5265_), .Y(_5266_) );
	NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_4820_), .B(_4926_), .Y(_5267_) );
	XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(_4822_), .Y(_5268_) );
	INVX1 INVX1_869 ( .gnd(gnd), .vdd(vdd), .A(_5268_), .Y(_5269_) );
	NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_5269_), .B(divider_divuResult_10_bF_buf1), .Y(_5270_) );
	NAND3X1 NAND3X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .B(_4819_), .C(_4937__bF_buf0), .Y(_5271_) );
	NAND3X1 NAND3X1_1117 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .B(_5271_), .C(_5270_), .Y(_5272_) );
	NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_5268_), .B(divider_divuResult_10_bF_buf0), .Y(_5273_) );
	NAND3X1 NAND3X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_4923_), .B(_4924_), .C(_4937__bF_buf5), .Y(_5275_) );
	NAND3X1 NAND3X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_5275_), .C(_5273_), .Y(_5276_) );
	NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_5272_), .B(_5276_), .Y(_5277_) );
	INVX1 INVX1_870 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_9_), .Y(_5278_) );
	INVX1 INVX1_871 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_8_), .Y(_5279_) );
	NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf0), .B(_5279_), .Y(_5280_) );
	INVX1 INVX1_872 ( .gnd(gnd), .vdd(vdd), .A(_5280_), .Y(_5281_) );
	NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_8_), .B(_1746__bF_buf0), .Y(_5282_) );
	OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(_5282_), .C(_5281_), .Y(_5283_) );
	NAND3X1 NAND3X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_5283_), .B(_5266_), .C(_5277_), .Y(_5284_) );
	OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_4937__bF_buf4), .B(_5268_), .C(_5271_), .Y(_5286_) );
	INVX1 INVX1_873 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .Y(_5287_) );
	OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_5286_), .C(_5260_), .Y(_5288_) );
	OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_5287_), .C(_5288_), .Y(_5289_) );
	AOI21X1 AOI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_5284_), .B(_5289_), .C(_5254_), .Y(_5290_) );
	NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .B(_5278_), .Y(_5291_) );
	NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_9_), .B(_1746__bF_buf5), .Y(_5292_) );
	NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_5291_), .B(_5292_), .Y(_5293_) );
	INVX1 INVX1_874 ( .gnd(gnd), .vdd(vdd), .A(_5293_), .Y(_5294_) );
	NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_8_), .B(_5294_), .Y(_5295_) );
	NAND3X1 NAND3X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .B(_5266_), .C(_5277_), .Y(_5297_) );
	NAND3X1 NAND3X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf5), .B(_5235_), .C(_5237_), .Y(_5298_) );
	AOI21X1 AOI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_5237_), .B(_5235_), .C(_1735__bF_buf4), .Y(_5299_) );
	NAND3X1 NAND3X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf7), .B(_5245_), .C(_5246_), .Y(_5300_) );
	AOI21X1 AOI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_5298_), .B(_5300_), .C(_5299_), .Y(_5301_) );
	NAND3X1 NAND3X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_5210_), .C(_5202_), .Y(_5302_) );
	AOI21X1 AOI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_5202_), .B(_5210_), .C(_4999__bF_buf0), .Y(_5303_) );
	NAND3X1 NAND3X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf6), .B(_5221_), .C(_5223_), .Y(_5304_) );
	OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_5304_), .B(_5303_), .C(_5302_), .Y(_5305_) );
	AOI21X1 AOI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_5229_), .B(_5301_), .C(_5305_), .Y(_5306_) );
	OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_5254_), .B(_5297_), .C(_5306_), .Y(_5308_) );
	NAND3X1 NAND3X1_1126 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .B(_5148_), .C(_5154_), .Y(_5309_) );
	NAND3X1 NAND3X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf4), .B(_5157_), .C(_5160_), .Y(_5310_) );
	NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_5309_), .B(_5310_), .Y(_5311_) );
	INVX1 INVX1_875 ( .gnd(gnd), .vdd(vdd), .A(_5195_), .Y(_5312_) );
	NAND3X1 NAND3X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf1), .B(_5312_), .C(_5126__bF_buf3), .Y(_5313_) );
	NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_4937__bF_buf3), .Y(_5314_) );
	NAND3X1 NAND3X1_1129 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .B(_5313_), .C(_5314_), .Y(_5315_) );
	NAND3X1 NAND3X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf3), .B(_5196_), .C(_5194_), .Y(_5316_) );
	NAND3X1 NAND3X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_4748_), .B(_4867_), .C(_4937__bF_buf2), .Y(_5317_) );
	NAND3X1 NAND3X1_1132 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .B(_5188_), .C(_5317_), .Y(_5319_) );
	NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_4759_), .B(_4937__bF_buf1), .Y(_5320_) );
	XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_5185_), .B(_5180_), .Y(_5321_) );
	NAND3X1 NAND3X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_3171__bF_buf0), .B(_5126__bF_buf2), .C(_5321_), .Y(_5322_) );
	NAND3X1 NAND3X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf0), .B(_5322_), .C(_5320_), .Y(_5323_) );
	AOI22X1 AOI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_5315_), .B(_5316_), .C(_5319_), .D(_5323_), .Y(_5324_) );
	NAND3X1 NAND3X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_5176_), .B(_5324_), .C(_5311_), .Y(_5325_) );
	NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_5146_), .B(_5325_), .C(_5112_), .Y(_5326_) );
	OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(_5308_), .C(_5326_), .Y(_5327_) );
	NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_5327_), .Y(_5328_) );
	NAND3X1 NAND3X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_5069_), .C(_5328_), .Y(_5330_) );
	AOI21X1 AOI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_5330_), .B(_5058_), .C(_3260_), .Y(divider_divuResult_9_) );
	OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf5), .B(_4938_), .Y(_5331_) );
	INVX8 INVX8_37 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .Y(_5332_) );
	NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(divider_divuResult_9_bF_buf4), .Y(_5333_) );
	OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf3), .B(_5333_), .C(divider_absoluteValue_B_flipSign_result_23_bF_buf1), .Y(_5334_) );
	OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(divider_divuResult_9_bF_buf3), .C(_2229__bF_buf1), .Y(_5335_) );
	OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_5335_), .B(divider_absoluteValue_B_flipSign_result_23_bF_buf0), .Y(_5336_) );
	NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_4956_), .B(_4950_), .Y(_5337_) );
	INVX1 INVX1_876 ( .gnd(gnd), .vdd(vdd), .A(_4986_), .Y(_5338_) );
	INVX1 INVX1_877 ( .gnd(gnd), .vdd(vdd), .A(_5069_), .Y(_5340_) );
	AOI21X1 AOI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_5327_), .B(_5201_), .C(_5340_), .Y(_5341_) );
	OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_5049_), .B(_5341_), .C(_5338_), .Y(_5342_) );
	AOI21X1 AOI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_5342_), .B(_5052_), .C(_5337_), .Y(_5343_) );
	NAND3X1 NAND3X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_5337_), .B(_5052_), .C(_5342_), .Y(_5344_) );
	INVX1 INVX1_878 ( .gnd(gnd), .vdd(vdd), .A(_5344_), .Y(_5345_) );
	OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .B(_5345_), .C(divider_divuResult_9_bF_buf2), .Y(_5346_) );
	OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_4948_), .B(divider_divuResult_10_bF_buf5), .C(_4947_), .Y(_5347_) );
	NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_5069_), .B(_4987_), .Y(_5348_) );
	OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_5348_), .C(_5058_), .Y(_5349_) );
	AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_5253_), .B(_5229_), .Y(_5351_) );
	NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_5289_), .B(_5284_), .Y(_5352_) );
	NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_5351_), .B(_5352_), .Y(_5353_) );
	NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_5260_), .B(_5265_), .Y(_5354_) );
	NAND3X1 NAND3X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_5271_), .C(_5270_), .Y(_5355_) );
	NAND3X1 NAND3X1_1139 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_5275_), .C(_5273_), .Y(_5356_) );
	NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_5355_), .B(_5356_), .Y(_5357_) );
	INVX1 INVX1_879 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .Y(_5358_) );
	NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_5358_), .C(_5357_), .Y(_5359_) );
	NOR3X1 NOR3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf6), .B(_5213_), .C(_5214_), .Y(_5360_) );
	AOI21X1 AOI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_5202_), .B(_5210_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .Y(_5362_) );
	NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_5224_), .B(_5228_), .Y(_5363_) );
	OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_5362_), .B(_5360_), .C(_5363_), .Y(_5364_) );
	OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_5240_), .B(_5239_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .Y(_5365_) );
	NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_5298_), .B(_5300_), .Y(_5366_) );
	NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .B(_5366_), .Y(_5367_) );
	INVX1 INVX1_880 ( .gnd(gnd), .vdd(vdd), .A(_5302_), .Y(_5368_) );
	OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_5213_), .B(_5214_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .Y(_5369_) );
	INVX1 INVX1_881 ( .gnd(gnd), .vdd(vdd), .A(_5304_), .Y(_5370_) );
	AOI21X1 AOI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_5370_), .B(_5369_), .C(_5368_), .Y(_5371_) );
	OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_5367_), .B(_5364_), .C(_5371_), .Y(_5373_) );
	AOI21X1 AOI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_5351_), .B(_5359_), .C(_5373_), .Y(_5374_) );
	NAND3X1 NAND3X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_5326_), .B(_5069_), .C(_4987_), .Y(_5375_) );
	AOI21X1 AOI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_5353_), .B(_5374_), .C(_5375_), .Y(_5376_) );
	OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_5376_), .B(_5349_), .C(_3261__bF_buf2), .Y(_5377_) );
	NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_5347_), .B(_5377__bF_buf5), .Y(_5378_) );
	NAND3X1 NAND3X1_1141 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf3), .B(_5378_), .C(_5346_), .Y(_5379_) );
	INVX1 INVX1_882 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .Y(_5380_) );
	NAND3X1 NAND3X1_1142 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf1), .B(_5344_), .C(_5380_), .Y(_5381_) );
	INVX1 INVX1_883 ( .gnd(gnd), .vdd(vdd), .A(_5347_), .Y(_5382_) );
	NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_5382_), .B(_5377__bF_buf4), .Y(_5384_) );
	NAND3X1 NAND3X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf2), .B(_5384_), .C(_5381_), .Y(_5385_) );
	AOI22X1 AOI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_5334_), .B(_5336_), .C(_5379_), .D(_5385_), .Y(_5386_) );
	OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_4959_), .B(_4973_), .C(_5377__bF_buf3), .Y(_5387_) );
	INVX1 INVX1_884 ( .gnd(gnd), .vdd(vdd), .A(_4974_), .Y(_5388_) );
	NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_5050_), .B(_5388_), .Y(_5389_) );
	OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_5049_), .B(_5341_), .C(_4985_), .Y(_5390_) );
	NAND3X1 NAND3X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_5389_), .B(_4980_), .C(_5390_), .Y(_5391_) );
	INVX1 INVX1_885 ( .gnd(gnd), .vdd(vdd), .A(_5389_), .Y(_5392_) );
	OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_4978_), .B(divider_divuResult_10_bF_buf4), .C(_4983_), .Y(_5393_) );
	INVX1 INVX1_886 ( .gnd(gnd), .vdd(vdd), .A(_5393_), .Y(_5395_) );
	NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf3), .B(_5395_), .Y(_5396_) );
	INVX1 INVX1_887 ( .gnd(gnd), .vdd(vdd), .A(_5396_), .Y(_5397_) );
	NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf3), .B(_5393_), .Y(_5398_) );
	INVX1 INVX1_888 ( .gnd(gnd), .vdd(vdd), .A(_5398_), .Y(_5399_) );
	INVX1 INVX1_889 ( .gnd(gnd), .vdd(vdd), .A(_5049_), .Y(_5400_) );
	AOI21X1 AOI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_5103_), .B(_5100_), .C(_1505__bF_buf4), .Y(_5401_) );
	OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .B(_5107_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .Y(_5402_) );
	NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .B(_5402_), .Y(_5403_) );
	NOR3X1 NOR3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_5403_), .B(_5401_), .C(_5091_), .Y(_5404_) );
	INVX1 INVX1_890 ( .gnd(gnd), .vdd(vdd), .A(_5134_), .Y(_5406_) );
	NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .B(_5404_), .Y(_5407_) );
	INVX1 INVX1_891 ( .gnd(gnd), .vdd(vdd), .A(_5146_), .Y(_5408_) );
	NAND3X1 NAND3X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_5408_), .B(_5200_), .C(_5404_), .Y(_5409_) );
	NAND3X1 NAND3X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .B(_5407_), .C(_5409_), .Y(_5410_) );
	INVX1 INVX1_892 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .Y(_5411_) );
	NAND3X1 NAND3X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_5408_), .B(_5411_), .C(_5404_), .Y(_5412_) );
	AOI21X1 AOI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_5353_), .B(_5374_), .C(_5412_), .Y(_5413_) );
	OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_5410_), .B(_5413_), .C(_5069_), .Y(_5414_) );
	AOI22X1 AOI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_5397_), .B(_5399_), .C(_5400_), .D(_5414_), .Y(_5415_) );
	OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_5415_), .C(_5392_), .Y(_5417_) );
	NAND3X1 NAND3X1_1148 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf0), .B(_5391_), .C(_5417_), .Y(_5418_) );
	NAND3X1 NAND3X1_1149 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf1), .B(_5387_), .C(_5418_), .Y(_5419_) );
	INVX1 INVX1_893 ( .gnd(gnd), .vdd(vdd), .A(_5387_), .Y(_5420_) );
	OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_5415_), .C(_5389_), .Y(_5421_) );
	NAND3X1 NAND3X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_5392_), .B(_4980_), .C(_5390_), .Y(_5422_) );
	AOI21X1 AOI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_5421_), .B(_5422_), .C(_5377__bF_buf2), .Y(_5423_) );
	OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .B(_5423_), .C(_4424__bF_buf1), .Y(_5424_) );
	NOR3X1 NOR3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_4985_), .B(_5049_), .C(_5341_), .Y(_5425_) );
	OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_5415_), .B(_5425_), .C(divider_divuResult_9_bF_buf5), .Y(_5426_) );
	NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_5395_), .B(_5377__bF_buf1), .Y(_5427_) );
	NAND3X1 NAND3X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf3), .B(_5427_), .C(_5426_), .Y(_5428_) );
	INVX1 INVX1_894 ( .gnd(gnd), .vdd(vdd), .A(_4985_), .Y(_5429_) );
	NAND3X1 NAND3X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_5429_), .B(_5400_), .C(_5414_), .Y(_5430_) );
	AOI21X1 AOI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_5390_), .B(_5430_), .C(_5377__bF_buf0), .Y(_5431_) );
	NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_5393_), .B(divider_divuResult_9_bF_buf4), .Y(_5432_) );
	OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_5431_), .B(_5432_), .C(divider_absoluteValue_B_flipSign_result_20_bF_buf2), .Y(_5433_) );
	NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_5428_), .B(_5433_), .Y(_5434_) );
	AOI21X1 AOI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_5424_), .B(_5419_), .C(_5434_), .Y(_5435_) );
	NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(_5435_), .Y(_5436_) );
	NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_4989_), .B(_5003_), .Y(_5439_) );
	OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf3), .B(_5439_), .Y(_5440_) );
	INVX1 INVX1_895 ( .gnd(gnd), .vdd(vdd), .A(_5011_), .Y(_5441_) );
	NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_5441_), .B(_5005_), .Y(_5442_) );
	INVX1 INVX1_896 ( .gnd(gnd), .vdd(vdd), .A(_5048_), .Y(_5443_) );
	AOI21X1 AOI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_5327_), .B(_5201_), .C(_5068_), .Y(_5444_) );
	OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_5443_), .B(_5444_), .C(_5023_), .Y(_5445_) );
	NAND3X1 NAND3X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_5017_), .B(_5442_), .C(_5445_), .Y(_5446_) );
	INVX1 INVX1_897 ( .gnd(gnd), .vdd(vdd), .A(_5017_), .Y(_5447_) );
	INVX1 INVX1_898 ( .gnd(gnd), .vdd(vdd), .A(_5442_), .Y(_5448_) );
	INVX1 INVX1_899 ( .gnd(gnd), .vdd(vdd), .A(_5068_), .Y(_5450_) );
	OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_5410_), .B(_5413_), .C(_5450_), .Y(_5451_) );
	AOI22X1 AOI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(_5022_), .C(_5048_), .D(_5451_), .Y(_5452_) );
	OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_5447_), .B(_5452_), .C(_5448_), .Y(_5453_) );
	NAND3X1 NAND3X1_1154 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf2), .B(_5446_), .C(_5453_), .Y(_5454_) );
	NAND3X1 NAND3X1_1155 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf2), .B(_5440_), .C(_5454_), .Y(_5455_) );
	NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_5439_), .B(_5377__bF_buf5), .Y(_5456_) );
	OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_5447_), .B(_5452_), .C(_5442_), .Y(_5457_) );
	NAND3X1 NAND3X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_5017_), .B(_5448_), .C(_5445_), .Y(_5458_) );
	NAND3X1 NAND3X1_1157 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf1), .B(_5458_), .C(_5457_), .Y(_5459_) );
	NAND3X1 NAND3X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf2), .B(_5456_), .C(_5459_), .Y(_5461_) );
	INVX1 INVX1_900 ( .gnd(gnd), .vdd(vdd), .A(_5023_), .Y(_5462_) );
	NAND3X1 NAND3X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_5462_), .B(_5048_), .C(_5451_), .Y(_5463_) );
	AOI21X1 AOI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_5445_), .B(_5463_), .C(_5377__bF_buf4), .Y(_5464_) );
	INVX1 INVX1_901 ( .gnd(gnd), .vdd(vdd), .A(_5464_), .Y(_5465_) );
	OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf0), .B(_5016_), .Y(_5466_) );
	NAND3X1 NAND3X1_1160 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf0), .B(_5466_), .C(_5465_), .Y(_5467_) );
	NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(divider_divuResult_9_bF_buf5), .Y(_5468_) );
	OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_5464_), .B(_5468_), .C(_3263__bF_buf0), .Y(_5469_) );
	AOI22X1 AOI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_5467_), .B(_5469_), .C(_5455_), .D(_5461_), .Y(_5470_) );
	OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_4599_), .B(divider_divuResult_10_bF_buf3), .C(_5063_), .Y(_5472_) );
	INVX1 INVX1_902 ( .gnd(gnd), .vdd(vdd), .A(_5472_), .Y(_5473_) );
	NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_5473_), .B(divider_divuResult_9_bF_buf4), .Y(_5474_) );
	NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_5059_), .B(_5064_), .Y(_5475_) );
	INVX1 INVX1_903 ( .gnd(gnd), .vdd(vdd), .A(_5475_), .Y(_5476_) );
	NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .B(_5066_), .Y(_5477_) );
	AOI21X1 AOI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_5327_), .B(_5201_), .C(_5477_), .Y(_5478_) );
	OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(_5478_), .C(_5476_), .Y(_5479_) );
	INVX1 INVX1_904 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .Y(_5480_) );
	OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_5066_), .B(_5067_), .C(_5328_), .Y(_5481_) );
	NAND3X1 NAND3X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_5480_), .B(_5475_), .C(_5481_), .Y(_5483_) );
	AOI21X1 AOI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_5483_), .B(_5479_), .C(_5377__bF_buf3), .Y(_5484_) );
	OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_5484_), .B(_5474_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .Y(_5485_) );
	NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_5472_), .B(_5377__bF_buf2), .Y(_5486_) );
	NAND3X1 NAND3X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_5480_), .B(_5476_), .C(_5481_), .Y(_5487_) );
	OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(_5478_), .C(_5475_), .Y(_5488_) );
	NAND3X1 NAND3X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_5487_), .B(_5488_), .C(divider_divuResult_9_bF_buf3), .Y(_5489_) );
	NAND3X1 NAND3X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf1), .B(_5486_), .C(_5489_), .Y(_5490_) );
	INVX1 INVX1_905 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .Y(_5491_) );
	AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_4987_), .B(_5069_), .Y(_5492_) );
	NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_5410_), .B(_5492_), .Y(_5494_) );
	AOI21X1 AOI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_5272_), .B(_5276_), .C(_5354_), .Y(_5495_) );
	AOI22X1 AOI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_5356_), .B(_5288_), .C(_5283_), .D(_5495_), .Y(_5496_) );
	OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_5254_), .B(_5496_), .C(_5374_), .Y(_5497_) );
	NAND3X1 NAND3X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_5497_), .B(_5326_), .C(_5492_), .Y(_5498_) );
	NAND3X1 NAND3X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_5058_), .B(_5494_), .C(_5498_), .Y(_5499_) );
	NAND3X1 NAND3X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_5477_), .B(_5201_), .C(_5327_), .Y(_5500_) );
	NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_5500_), .B(_5481_), .Y(_5501_) );
	NAND3X1 NAND3X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf1), .B(_5499__bF_buf3), .C(_5501_), .Y(_5502_) );
	OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_5491_), .B(divider_divuResult_9_bF_buf2), .C(_5502_), .Y(_5503_) );
	OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf4), .B(_5503_), .C(_5490_), .Y(_5505_) );
	AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_5505_), .B(_5485_), .Y(_5506_) );
	NAND3X1 NAND3X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf1), .B(_5440_), .C(_5454_), .Y(_5507_) );
	AOI21X1 AOI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_5454_), .B(_5440_), .C(_3789__bF_buf0), .Y(_5508_) );
	NAND3X1 NAND3X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf3), .B(_5466_), .C(_5465_), .Y(_5509_) );
	OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_5509_), .B(_5508_), .C(_5507_), .Y(_5510_) );
	AOI21X1 AOI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_5506_), .B(_5470_), .C(_5510_), .Y(_5511_) );
	NAND3X1 NAND3X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf0), .B(_5387_), .C(_5418_), .Y(_5512_) );
	AOI21X1 AOI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_5418_), .B(_5387_), .C(_4424__bF_buf3), .Y(_5513_) );
	AOI21X1 AOI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_5512_), .B(_5428_), .C(_5513_), .Y(_5514_) );
	INVX8 INVX8_38 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf3), .Y(_5516_) );
	OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf2), .B(_5333_), .C(_5516__bF_buf3), .Y(_5517_) );
	NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf2), .B(_5335_), .Y(_5518_) );
	NAND3X1 NAND3X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf1), .B(_5378_), .C(_5346_), .Y(_5519_) );
	OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_5518_), .B(_5519_), .C(_5517_), .Y(_5520_) );
	AOI21X1 AOI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(_5514_), .C(_5520_), .Y(_5521_) );
	OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_5436_), .B(_5511_), .C(_5521_), .Y(_5522_) );
	NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_5334_), .B(_5336_), .Y(_5523_) );
	NAND3X1 NAND3X1_1173 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf2), .B(_5384_), .C(_5381_), .Y(_5524_) );
	NAND3X1 NAND3X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_5519_), .B(_5524_), .C(_5523_), .Y(_5525_) );
	OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .B(_5423_), .C(divider_absoluteValue_B_flipSign_result_21_bF_buf0), .Y(_5527_) );
	AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_5433_), .B(_5428_), .Y(_5528_) );
	NAND3X1 NAND3X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_5512_), .B(_5527_), .C(_5528_), .Y(_5529_) );
	NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_5455_), .B(_5461_), .Y(_5530_) );
	NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_5469_), .B(_5467_), .Y(_5531_) );
	NAND3X1 NAND3X1_1176 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .B(_5486_), .C(_5489_), .Y(_5532_) );
	OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_5484_), .B(_5474_), .C(_2887__bF_buf0), .Y(_5533_) );
	NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_5377__bF_buf1), .Y(_5534_) );
	NAND3X1 NAND3X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf1), .B(_5502_), .C(_5534_), .Y(_5535_) );
	NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_5491_), .B(_5377__bF_buf0), .Y(_5536_) );
	INVX1 INVX1_906 ( .gnd(gnd), .vdd(vdd), .A(_5500_), .Y(_5538_) );
	NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_5478_), .B(_5538_), .Y(_5539_) );
	NAND3X1 NAND3X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf0), .B(_5499__bF_buf2), .C(_5539_), .Y(_5540_) );
	NAND3X1 NAND3X1_1179 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf3), .B(_5536_), .C(_5540_), .Y(_5541_) );
	NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_5535_), .B(_5541_), .Y(_5542_) );
	AOI21X1 AOI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_5532_), .B(_5533_), .C(_5542_), .Y(_5543_) );
	NAND3X1 NAND3X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_5531_), .B(_5543_), .C(_5530_), .Y(_5544_) );
	NOR3X1 NOR3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_5525_), .B(_5529_), .C(_5544_), .Y(_5545_) );
	OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_5071_), .B(divider_divuResult_10_bF_buf2), .C(_5103_), .Y(_5546_) );
	NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_5377__bF_buf5), .Y(_5547_) );
	NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_5401_), .B(_5091_), .Y(_5549_) );
	INVX1 INVX1_907 ( .gnd(gnd), .vdd(vdd), .A(_5200_), .Y(_5550_) );
	OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(_5308_), .C(_5411_), .Y(_5551_) );
	AOI21X1 AOI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_5551_), .B(_5550_), .C(_5146_), .Y(_5552_) );
	OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .B(_5552_), .C(_5111_), .Y(_5553_) );
	NAND3X1 NAND3X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .B(_5549_), .C(_5553_), .Y(_5554_) );
	INVX1 INVX1_908 ( .gnd(gnd), .vdd(vdd), .A(_5549_), .Y(_5555_) );
	AOI21X1 AOI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_5374_), .B(_5353_), .C(_5325_), .Y(_5556_) );
	OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_5200_), .B(_5556_), .C(_5408_), .Y(_5557_) );
	AOI22X1 AOI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_5110_), .C(_5134_), .D(_5557_), .Y(_5558_) );
	OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .B(_5558_), .C(_5555_), .Y(_5560_) );
	NAND3X1 NAND3X1_1182 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf1), .B(_5554_), .C(_5560_), .Y(_5561_) );
	NAND3X1 NAND3X1_1183 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .B(_5547_), .C(_5561_), .Y(_5562_) );
	INVX1 INVX1_909 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .Y(_5563_) );
	NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_5563_), .B(_5377__bF_buf4), .Y(_5564_) );
	OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_5097_), .B(_5558_), .C(_5549_), .Y(_5565_) );
	NAND3X1 NAND3X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .B(_5555_), .C(_5553_), .Y(_5566_) );
	NAND3X1 NAND3X1_1185 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf0), .B(_5566_), .C(_5565_), .Y(_5567_) );
	NAND3X1 NAND3X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf2), .B(_5564_), .C(_5567_), .Y(_5568_) );
	NOR3X1 NOR3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_5111_), .B(_5406_), .C(_5552_), .Y(_5569_) );
	OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_5558_), .B(_5569_), .C(divider_divuResult_9_bF_buf5), .Y(_5571_) );
	OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_5108_), .C(_5377__bF_buf3), .Y(_5572_) );
	NAND3X1 NAND3X1_1187 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .B(_5572_), .C(_5571_), .Y(_5573_) );
	NAND3X1 NAND3X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_5403_), .B(_5134_), .C(_5557_), .Y(_5574_) );
	AOI21X1 AOI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_5553_), .B(_5574_), .C(_5377__bF_buf2), .Y(_5575_) );
	NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5094_), .Y(_5576_) );
	INVX1 INVX1_910 ( .gnd(gnd), .vdd(vdd), .A(_5576_), .Y(_5577_) );
	AOI21X1 AOI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_5499__bF_buf1), .B(_3261__bF_buf3), .C(_5577_), .Y(_5578_) );
	OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_5578_), .B(_5575_), .C(_1505__bF_buf3), .Y(_5579_) );
	AOI22X1 AOI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .B(_5579_), .C(_5562_), .D(_5568_), .Y(_5580_) );
	NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_5550_), .B(_5551_), .Y(_5582_) );
	XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_5582_), .B(_5145_), .Y(_5583_) );
	NAND3X1 NAND3X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf2), .B(_5499__bF_buf0), .C(_5583_), .Y(_5584_) );
	OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(divider_divuResult_10_bF_buf1), .C(_5129_), .Y(_5585_) );
	NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_5585_), .B(_5377__bF_buf1), .Y(_5586_) );
	NAND3X1 NAND3X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf0), .B(_5586_), .C(_5584_), .Y(_5587_) );
	INVX1 INVX1_911 ( .gnd(gnd), .vdd(vdd), .A(_5585_), .Y(_5588_) );
	NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_5588_), .B(_5377__bF_buf0), .Y(_5589_) );
	INVX1 INVX1_912 ( .gnd(gnd), .vdd(vdd), .A(_5145_), .Y(_5590_) );
	XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_5582_), .B(_5590_), .Y(_5591_) );
	NAND3X1 NAND3X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf1), .B(_5499__bF_buf3), .C(_5591_), .Y(_5593_) );
	NAND3X1 NAND3X1_1192 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .B(_5589_), .C(_5593_), .Y(_5594_) );
	NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_5594_), .Y(_5595_) );
	OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_5123_), .C(_5377__bF_buf5), .Y(_5596_) );
	OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5138_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .Y(_5597_) );
	OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .B(_5114_), .C(_1484__bF_buf4), .Y(_5598_) );
	NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_5598_), .B(_5597_), .Y(_5599_) );
	AOI21X1 AOI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_5551_), .B(_5550_), .C(_5590_), .Y(_5600_) );
	INVX1 INVX1_913 ( .gnd(gnd), .vdd(vdd), .A(_5600_), .Y(_5601_) );
	NAND3X1 NAND3X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_5599_), .C(_5601_), .Y(_5602_) );
	INVX1 INVX1_914 ( .gnd(gnd), .vdd(vdd), .A(_5599_), .Y(_5604_) );
	OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_5600_), .C(_5604_), .Y(_5605_) );
	NAND3X1 NAND3X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_5602_), .B(_5605_), .C(divider_divuResult_9_bF_buf4), .Y(_5606_) );
	NAND3X1 NAND3X1_1195 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_5596_), .C(_5606_), .Y(_5607_) );
	OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5138_), .C(_5377__bF_buf4), .Y(_5608_) );
	OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_5600_), .C(_5599_), .Y(_5609_) );
	NAND3X1 NAND3X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_5604_), .C(_5601_), .Y(_5610_) );
	NAND3X1 NAND3X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_5609_), .B(_5610_), .C(divider_divuResult_9_bF_buf3), .Y(_5611_) );
	NAND3X1 NAND3X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf0), .B(_5608_), .C(_5611_), .Y(_5612_) );
	AOI21X1 AOI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_5607_), .B(_5612_), .C(_5595_), .Y(_5613_) );
	NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_5613_), .B(_5580_), .Y(_5615_) );
	NAND3X1 NAND3X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_5157_), .B(_5160_), .C(_5377__bF_buf3), .Y(_5616_) );
	INVX1 INVX1_915 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .Y(_5617_) );
	INVX1 INVX1_916 ( .gnd(gnd), .vdd(vdd), .A(_5176_), .Y(_5618_) );
	OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(_5308_), .C(_5324_), .Y(_5619_) );
	AOI21X1 AOI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_5619_), .B(_5199_), .C(_5618_), .Y(_5620_) );
	INVX1 INVX1_917 ( .gnd(gnd), .vdd(vdd), .A(_5620_), .Y(_5621_) );
	NAND3X1 NAND3X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_5617_), .B(_5311_), .C(_5621_), .Y(_5622_) );
	INVX1 INVX1_918 ( .gnd(gnd), .vdd(vdd), .A(_5311_), .Y(_5623_) );
	OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5620_), .C(_5623_), .Y(_5624_) );
	NAND3X1 NAND3X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_5622_), .B(_5624_), .C(divider_divuResult_9_bF_buf2), .Y(_5626_) );
	NAND3X1 NAND3X1_1202 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .B(_5616_), .C(_5626_), .Y(_5627_) );
	NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_5159_), .Y(_5628_) );
	OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_4937__bF_buf0), .B(_5628_), .C(_5157_), .Y(_5629_) );
	NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_5629_), .B(_5377__bF_buf2), .Y(_5630_) );
	OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5620_), .C(_5311_), .Y(_5631_) );
	NAND3X1 NAND3X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_5617_), .B(_5623_), .C(_5621_), .Y(_5632_) );
	NAND3X1 NAND3X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_5631_), .B(_5632_), .C(divider_divuResult_9_bF_buf1), .Y(_5633_) );
	NAND3X1 NAND3X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf1), .B(_5630_), .C(_5633_), .Y(_5634_) );
	NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_5627_), .B(_5634_), .Y(_5635_) );
	NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_5199_), .B(_5619_), .Y(_5637_) );
	XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_5637_), .B(_5176_), .Y(_5638_) );
	NAND3X1 NAND3X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf0), .B(_5499__bF_buf2), .C(_5638_), .Y(_5639_) );
	NAND3X1 NAND3X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_5163_), .B(_5166_), .C(_5377__bF_buf1), .Y(_5640_) );
	NAND3X1 NAND3X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf3), .B(_5639_), .C(_5640_), .Y(_5641_) );
	XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_5637_), .B(_5618_), .Y(_5642_) );
	NAND3X1 NAND3X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf3), .B(_5499__bF_buf1), .C(_5642_), .Y(_5643_) );
	OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_5171_), .B(divider_divuResult_10_bF_buf0), .C(_5163_), .Y(_5644_) );
	NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_5644_), .B(_5377__bF_buf0), .Y(_5645_) );
	NAND3X1 NAND3X1_1210 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .B(_5645_), .C(_5643_), .Y(_5646_) );
	AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_5641_), .B(_5646_), .Y(_5648_) );
	OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(divider_divuResult_10_bF_buf5), .C(_5196_), .Y(_5649_) );
	INVX1 INVX1_919 ( .gnd(gnd), .vdd(vdd), .A(_5649_), .Y(_5650_) );
	NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_5315_), .B(_5316_), .Y(_5651_) );
	OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_5290_), .B(_5308_), .C(_5651_), .Y(_5652_) );
	OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_5650_), .C(_5652_), .Y(_5653_) );
	INVX1 INVX1_920 ( .gnd(gnd), .vdd(vdd), .A(_5190_), .Y(_5654_) );
	NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_5191_), .B(_5654_), .Y(_5655_) );
	INVX1 INVX1_921 ( .gnd(gnd), .vdd(vdd), .A(_5655_), .Y(_5656_) );
	NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_5656_), .B(_5653_), .Y(_5657_) );
	INVX1 INVX1_922 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .Y(_5659_) );
	NAND3X1 NAND3X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_5659_), .B(_5655_), .C(_5652_), .Y(_5660_) );
	NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_5660_), .B(_5657_), .Y(_5661_) );
	NAND3X1 NAND3X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf2), .B(_5499__bF_buf0), .C(_5661_), .Y(_5662_) );
	NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_5189_), .B(_5377__bF_buf5), .Y(_5663_) );
	AOI21X1 AOI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_5663_), .B(_5662_), .C(_8971__bF_buf2), .Y(_5664_) );
	NAND3X1 NAND3X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf1), .B(_5662_), .C(_5663_), .Y(_5665_) );
	XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_5497_), .B(_5651_), .Y(_5666_) );
	NAND3X1 NAND3X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf1), .B(_5666_), .C(_5499__bF_buf3), .Y(_5667_) );
	NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_5650_), .B(_5377__bF_buf4), .Y(_5668_) );
	NAND3X1 NAND3X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf5), .B(_5667_), .C(_5668_), .Y(_5670_) );
	AOI21X1 AOI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_5665_), .B(_5670_), .C(_5664_), .Y(_5671_) );
	NAND3X1 NAND3X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_5671_), .B(_5635_), .C(_5648_), .Y(_5672_) );
	OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_5629_), .B(divider_divuResult_9_bF_buf0), .C(_5626_), .Y(_5673_) );
	NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .B(_5673_), .Y(_5674_) );
	NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .B(_5673_), .Y(_5675_) );
	INVX1 INVX1_923 ( .gnd(gnd), .vdd(vdd), .A(_5641_), .Y(_5676_) );
	AOI21X1 AOI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_5676_), .B(_5675_), .C(_5674_), .Y(_5677_) );
	AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_5672_), .B(_5677_), .Y(_5678_) );
	NAND3X1 NAND3X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf1), .B(_5547_), .C(_5561_), .Y(_5679_) );
	AOI21X1 AOI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_5561_), .B(_5547_), .C(_1944__bF_buf0), .Y(_5681_) );
	OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_5577_), .B(divider_divuResult_9_bF_buf5), .C(_5571_), .Y(_5682_) );
	OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_5682_), .B(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .Y(_5683_) );
	OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_5681_), .B(_5683_), .C(_5679_), .Y(_5684_) );
	NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_5609_), .B(_5610_), .Y(_5685_) );
	OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_5377__bF_buf3), .B(_5685_), .C(_5608_), .Y(_5686_) );
	INVX1 INVX1_924 ( .gnd(gnd), .vdd(vdd), .A(_5686_), .Y(_5687_) );
	INVX1 INVX1_925 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .Y(_5688_) );
	OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf4), .B(_5686_), .C(_5688_), .Y(_5689_) );
	OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .B(_5687_), .C(_5689_), .Y(_5690_) );
	AOI21X1 AOI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_5690_), .B(_5580_), .C(_5684_), .Y(_5692_) );
	OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_5615_), .B(_5678_), .C(_5692_), .Y(_5693_) );
	AOI21X1 AOI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_5693_), .B(_5545_), .C(_5522_), .Y(_5694_) );
	NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_5215_), .Y(_5695_) );
	INVX1 INVX1_926 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .Y(_5696_) );
	NAND3X1 NAND3X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_5289_), .B(_5284_), .C(_5297_), .Y(_5697_) );
	AOI21X1 AOI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_5697_), .B(_5253_), .C(_5301_), .Y(_5698_) );
	OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_5696_), .B(_5698_), .C(_5304_), .Y(_5699_) );
	XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_5699_), .B(_5695_), .Y(_5700_) );
	OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_5213_), .B(_5214_), .C(_5377__bF_buf2), .Y(_5701_) );
	OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_5377__bF_buf1), .B(_5700_), .C(_5701_), .Y(_5703_) );
	NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(_5703_), .Y(_5704_) );
	XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_5699_), .B(_5695_), .Y(_5705_) );
	NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .B(divider_divuResult_9_bF_buf4), .Y(_5706_) );
	NAND3X1 NAND3X1_1219 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .B(_5701_), .C(_5706_), .Y(_5707_) );
	NAND3X1 NAND3X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf0), .B(_5499__bF_buf2), .C(_5700_), .Y(_5708_) );
	NAND3X1 NAND3X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_5202_), .B(_5210_), .C(_5377__bF_buf0), .Y(_5709_) );
	NAND3X1 NAND3X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf2), .B(_5708_), .C(_5709_), .Y(_5710_) );
	XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_5698_), .B(_5363_), .Y(_5711_) );
	INVX1 INVX1_927 ( .gnd(gnd), .vdd(vdd), .A(_5711_), .Y(_5712_) );
	NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_5712_), .B(divider_divuResult_9_bF_buf3), .Y(_5714_) );
	NAND3X1 NAND3X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_5225_), .B(_5227_), .C(_5377__bF_buf5), .Y(_5715_) );
	NAND3X1 NAND3X1_1224 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_5715_), .C(_5714_), .Y(_5716_) );
	NAND3X1 NAND3X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_5221_), .B(_5223_), .C(_5377__bF_buf4), .Y(_5717_) );
	NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_5711_), .B(divider_divuResult_9_bF_buf2), .Y(_5718_) );
	NAND3X1 NAND3X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_5717_), .C(_5718_), .Y(_5719_) );
	AOI22X1 AOI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_5707_), .B(_5710_), .C(_5716_), .D(_5719_), .Y(_5720_) );
	NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_5238_), .B(_5242_), .Y(_5721_) );
	INVX1 INVX1_928 ( .gnd(gnd), .vdd(vdd), .A(_5300_), .Y(_5722_) );
	AOI22X1 AOI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(_5247_), .B(_5251_), .C(_5297_), .D(_5496_), .Y(_5723_) );
	OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_5722_), .B(_5723_), .C(_5721_), .Y(_5725_) );
	NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_5722_), .B(_5723_), .Y(_5726_) );
	NAND3X1 NAND3X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_5238_), .B(_5242_), .C(_5726_), .Y(_5727_) );
	NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_5725_), .B(_5727_), .Y(_5728_) );
	NAND3X1 NAND3X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf3), .B(_5728_), .C(_5499__bF_buf1), .Y(_5729_) );
	OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_5239_), .B(_5240_), .C(_5377__bF_buf3), .Y(_5730_) );
	AOI21X1 AOI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_5730_), .B(_5729_), .C(_4100__bF_buf5), .Y(_5731_) );
	NAND3X1 NAND3X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf4), .B(_5729_), .C(_5730_), .Y(_5732_) );
	NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_5247_), .B(_5251_), .Y(_5733_) );
	NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_5733_), .B(_5697_), .Y(_5734_) );
	NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_5723_), .B(_5734_), .Y(_5736_) );
	INVX1 INVX1_929 ( .gnd(gnd), .vdd(vdd), .A(_5736_), .Y(_5737_) );
	NAND3X1 NAND3X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf2), .B(_5737_), .C(_5499__bF_buf0), .Y(_5738_) );
	OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_5249_), .B(divider_divuResult_10_bF_buf4), .C(_5245_), .Y(_5739_) );
	NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_5739_), .B(_5377__bF_buf2), .Y(_5740_) );
	NAND3X1 NAND3X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_5738_), .C(_5740_), .Y(_5741_) );
	AOI21X1 AOI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .B(_5741_), .C(_5731_), .Y(_5742_) );
	NAND3X1 NAND3X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_5715_), .C(_5714_), .Y(_5743_) );
	OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .B(_5703_), .C(_5743_), .Y(_5744_) );
	AOI22X1 AOI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5744_), .C(_5742_), .D(_5720_), .Y(_5745_) );
	NAND3X1 NAND3X1_1233 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .B(_5729_), .C(_5730_), .Y(_5747_) );
	AOI21X1 AOI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_5725_), .B(_5727_), .C(_5377__bF_buf1), .Y(_5748_) );
	NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_5240_), .B(_5239_), .Y(_5749_) );
	AOI21X1 AOI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_5499__bF_buf3), .B(_3261__bF_buf1), .C(_5749_), .Y(_5750_) );
	OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_5750_), .B(_5748_), .C(_4100__bF_buf3), .Y(_5751_) );
	NAND3X1 NAND3X1_1234 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .B(_5738_), .C(_5740_), .Y(_5752_) );
	NAND3X1 NAND3X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_5245_), .B(_5246_), .C(_5377__bF_buf0), .Y(_5753_) );
	NAND3X1 NAND3X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf0), .B(_5736_), .C(_5499__bF_buf2), .Y(_5754_) );
	NAND3X1 NAND3X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_5754_), .C(_5753_), .Y(_5755_) );
	AOI22X1 AOI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_5752_), .B(_5755_), .C(_5747_), .D(_5751_), .Y(_5756_) );
	NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_5756_), .B(_5720_), .Y(_5758_) );
	NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .B(_5377__bF_buf5), .Y(_5759_) );
	OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_5292_), .B(_5354_), .C(_5260_), .Y(_5760_) );
	XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_5760_), .B(_5357_), .Y(_5761_) );
	INVX1 INVX1_930 ( .gnd(gnd), .vdd(vdd), .A(_5761_), .Y(_5762_) );
	NAND3X1 NAND3X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf3), .B(_5762_), .C(_5499__bF_buf1), .Y(_5763_) );
	NAND3X1 NAND3X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_5763_), .C(_5759_), .Y(_5764_) );
	AOI21X1 AOI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .B(_5763_), .C(_2470__bF_buf5), .Y(_5765_) );
	XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_5292_), .Y(_5766_) );
	INVX1 INVX1_931 ( .gnd(gnd), .vdd(vdd), .A(_5766_), .Y(_5767_) );
	NAND3X1 NAND3X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf2), .B(_5767_), .C(_5499__bF_buf0), .Y(_5769_) );
	OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_10_), .B(divider_divuResult_10_bF_buf3), .C(_5258_), .Y(_5770_) );
	NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_5770_), .B(_5377__bF_buf4), .Y(_5771_) );
	NAND3X1 NAND3X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_5769_), .C(_5771_), .Y(_5772_) );
	OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_5772_), .B(_5765_), .C(_5764_), .Y(_5773_) );
	NAND3X1 NAND3X1_1242 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .B(_5763_), .C(_5759_), .Y(_5774_) );
	NAND3X1 NAND3X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf1), .B(_5761_), .C(_5499__bF_buf3), .Y(_5775_) );
	NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_5287_), .B(_5377__bF_buf3), .Y(_5776_) );
	NAND3X1 NAND3X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf4), .B(_5775_), .C(_5776_), .Y(_5777_) );
	NAND3X1 NAND3X1_1245 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_5769_), .C(_5771_), .Y(_5778_) );
	NAND3X1 NAND3X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf0), .B(_5766_), .C(_5499__bF_buf2), .Y(_5780_) );
	INVX1 INVX1_932 ( .gnd(gnd), .vdd(vdd), .A(_5770_), .Y(_5781_) );
	NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_5781_), .B(_5377__bF_buf2), .Y(_5782_) );
	NAND3X1 NAND3X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_5780_), .C(_5782_), .Y(_5783_) );
	AOI22X1 AOI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(_5774_), .B(_5777_), .C(_5778_), .D(_5783_), .Y(_5784_) );
	NAND3X1 NAND3X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf3), .B(_5293_), .C(_5499__bF_buf1), .Y(_5785_) );
	NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(_5377__bF_buf1), .Y(_5786_) );
	NAND3X1 NAND3X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_5785_), .C(_5786_), .Y(_5787_) );
	AOI21X1 AOI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_5786_), .B(_5785_), .C(_1768__bF_buf4), .Y(_5788_) );
	OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_5282_), .B(_5788_), .C(_5787_), .Y(_5789_) );
	AOI21X1 AOI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_5789_), .B(_5784_), .C(_5773_), .Y(_5791_) );
	OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_5758_), .B(_5791_), .C(_5745_), .Y(_5792_) );
	NAND3X1 NAND3X1_1250 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .B(_5564_), .C(_5567_), .Y(_5793_) );
	NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .B(_5579_), .Y(_5794_) );
	NAND3X1 NAND3X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_5679_), .B(_5793_), .C(_5794_), .Y(_5795_) );
	AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_5594_), .Y(_5796_) );
	NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_5607_), .B(_5612_), .Y(_5797_) );
	NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_5797_), .B(_5796_), .Y(_5798_) );
	NAND3X1 NAND3X1_1252 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .B(_5662_), .C(_5663_), .Y(_5799_) );
	AOI21X1 AOI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_5657_), .B(_5660_), .C(_5377__bF_buf0), .Y(_5800_) );
	AOI22X1 AOI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_5317_), .B(_5188_), .C(_3261__bF_buf2), .D(_5499__bF_buf0), .Y(_5802_) );
	OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_5802_), .B(_5800_), .C(_8971__bF_buf0), .Y(_5803_) );
	NAND3X1 NAND3X1_1253 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .B(_5667_), .C(_5668_), .Y(_5804_) );
	INVX1 INVX1_933 ( .gnd(gnd), .vdd(vdd), .A(_5666_), .Y(_5805_) );
	NAND3X1 NAND3X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_3261__bF_buf1), .B(_5499__bF_buf3), .C(_5805_), .Y(_5806_) );
	NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_5649_), .B(_5377__bF_buf5), .Y(_5807_) );
	NAND3X1 NAND3X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf4), .B(_5806_), .C(_5807_), .Y(_5808_) );
	AOI22X1 AOI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_5804_), .B(_5808_), .C(_5799_), .D(_5803_), .Y(_5809_) );
	NAND3X1 NAND3X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .B(_5648_), .C(_5809_), .Y(_5810_) );
	NOR3X1 NOR3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_5798_), .B(_5795_), .C(_5810_), .Y(_5811_) );
	NAND3X1 NAND3X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_5792_), .B(_5811_), .C(_5545_), .Y(_5813_) );
	AOI21X1 AOI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_5694_), .B(_5813_), .C(_5332__bF_buf3), .Y(divider_divuResult_8_) );
	OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_5331_), .B(divider_divuResult_8_bF_buf6), .C(_2229__bF_buf0), .Y(_5814_) );
	XNOR2X1 XNOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_5814_), .B(divider_absoluteValue_B_flipSign_result_24_bF_buf1), .Y(_5815_) );
	NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_5379_), .B(_5385_), .Y(_5816_) );
	INVX1 INVX1_934 ( .gnd(gnd), .vdd(vdd), .A(_5816_), .Y(_5817_) );
	INVX1 INVX1_935 ( .gnd(gnd), .vdd(vdd), .A(_5512_), .Y(_5818_) );
	INVX1 INVX1_936 ( .gnd(gnd), .vdd(vdd), .A(_5428_), .Y(_5819_) );
	OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5818_), .C(_5527_), .Y(_5820_) );
	NAND3X1 NAND3X1_1258 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf1), .B(_5456_), .C(_5459_), .Y(_5821_) );
	NAND3X1 NAND3X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .B(_5821_), .C(_5531_), .Y(_5823_) );
	NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_5485_), .B(_5505_), .Y(_5824_) );
	INVX1 INVX1_937 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .Y(_5825_) );
	INVX1 INVX1_938 ( .gnd(gnd), .vdd(vdd), .A(_5509_), .Y(_5826_) );
	AOI21X1 AOI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_5821_), .B(_5826_), .C(_5825_), .Y(_5827_) );
	OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_5824_), .B(_5823_), .C(_5827_), .Y(_5828_) );
	NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_5798_), .B(_5795_), .Y(_5829_) );
	NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_5677_), .B(_5672_), .Y(_5830_) );
	AOI21X1 AOI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_5567_), .B(_5564_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .Y(_5831_) );
	NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf2), .B(_5682_), .Y(_5832_) );
	AOI21X1 AOI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_5832_), .B(_5793_), .C(_5831_), .Y(_5834_) );
	AOI21X1 AOI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_5611_), .B(_5608_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .Y(_5835_) );
	NAND3X1 NAND3X1_1260 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .B(_5608_), .C(_5611_), .Y(_5836_) );
	AOI21X1 AOI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_5688_), .B(_5836_), .C(_5835_), .Y(_5837_) );
	OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_5837_), .B(_5795_), .C(_5834_), .Y(_5838_) );
	AOI21X1 AOI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_5829_), .B(_5830_), .C(_5838_), .Y(_5839_) );
	NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_5792_), .B(_5811_), .Y(_5840_) );
	AOI21X1 AOI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_5840_), .B(_5839_), .C(_5544_), .Y(_5841_) );
	OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_5828_), .B(_5841_), .C(_5435_), .Y(_5842_) );
	AOI21X1 AOI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_5842_), .B(_5820_), .C(_5817_), .Y(_5843_) );
	NAND3X1 NAND3X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_5817_), .B(_5820_), .C(_5842_), .Y(_5845_) );
	INVX1 INVX1_939 ( .gnd(gnd), .vdd(vdd), .A(_5845_), .Y(_5846_) );
	OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_5843_), .B(_5846_), .C(divider_divuResult_8_bF_buf5), .Y(_5847_) );
	OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_5382_), .B(divider_divuResult_9_bF_buf1), .C(_5346_), .Y(_5848_) );
	AOI21X1 AOI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_5709_), .B(_5708_), .C(_4714__bF_buf1), .Y(_5849_) );
	AOI21X1 AOI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_5706_), .B(_5701_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .Y(_5850_) );
	AOI21X1 AOI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_5718_), .B(_5717_), .C(_4999__bF_buf3), .Y(_5851_) );
	AOI21X1 AOI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_5714_), .B(_5715_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .Y(_5852_) );
	OAI22X1 OAI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .B(_5850_), .C(_5851_), .D(_5852_), .Y(_5853_) );
	OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_5749_), .B(divider_divuResult_9_bF_buf0), .C(_5729_), .Y(_5854_) );
	INVX1 INVX1_940 ( .gnd(gnd), .vdd(vdd), .A(_5854_), .Y(_5856_) );
	OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .B(_5854_), .C(_5741_), .Y(_5857_) );
	OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_5856_), .C(_5857_), .Y(_5858_) );
	INVX1 INVX1_941 ( .gnd(gnd), .vdd(vdd), .A(_5703_), .Y(_5859_) );
	OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf0), .B(_5859_), .C(_5744_), .Y(_5860_) );
	OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_5853_), .B(_5858_), .C(_5860_), .Y(_5861_) );
	AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_5720_), .B(_5756_), .Y(_5862_) );
	INVX1 INVX1_942 ( .gnd(gnd), .vdd(vdd), .A(_5764_), .Y(_5863_) );
	OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_5287_), .B(divider_divuResult_9_bF_buf5), .C(_5763_), .Y(_5864_) );
	NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_5864_), .Y(_5865_) );
	AOI21X1 AOI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_5782_), .B(_5780_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .Y(_5867_) );
	AOI21X1 AOI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_5865_), .B(_5867_), .C(_5863_), .Y(_5868_) );
	AOI21X1 AOI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_5776_), .B(_5775_), .C(_2470__bF_buf3), .Y(_5869_) );
	AOI21X1 AOI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .B(_5763_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .Y(_5870_) );
	AOI21X1 AOI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_5782_), .B(_5780_), .C(_2547__bF_buf6), .Y(_5871_) );
	AOI21X1 AOI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_5771_), .B(_5769_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .Y(_5872_) );
	OAI22X1 OAI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_5869_), .B(_5870_), .C(_5871_), .D(_5872_), .Y(_5873_) );
	INVX1 INVX1_943 ( .gnd(gnd), .vdd(vdd), .A(_5282_), .Y(_5874_) );
	NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_9_), .B(_5377__bF_buf4), .Y(_5875_) );
	OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_5291_), .B(_5292_), .C(divider_divuResult_9_bF_buf4), .Y(_5876_) );
	AOI21X1 AOI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_5876_), .B(_5875_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .Y(_5878_) );
	NAND3X1 NAND3X1_1262 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .B(_5875_), .C(_5876_), .Y(_5879_) );
	AOI21X1 AOI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_5874_), .B(_5879_), .C(_5878_), .Y(_5880_) );
	OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_5873_), .B(_5880_), .C(_5868_), .Y(_5881_) );
	AOI21X1 AOI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_5862_), .B(_5881_), .C(_5861_), .Y(_5882_) );
	INVX1 INVX1_944 ( .gnd(gnd), .vdd(vdd), .A(_5810_), .Y(_5883_) );
	NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_5883_), .B(_5829_), .Y(_5884_) );
	OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_5882_), .B(_5884_), .C(_5839_), .Y(_5885_) );
	AOI21X1 AOI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_5885_), .B(_5545_), .C(_5522_), .Y(_5886_) );
	OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf2), .B(_5886__bF_buf3), .C(_5848_), .Y(_5887_) );
	NAND3X1 NAND3X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf1), .B(_5887_), .C(_5847_), .Y(_5889_) );
	INVX1 INVX1_945 ( .gnd(gnd), .vdd(vdd), .A(_5544_), .Y(_5890_) );
	AOI21X1 AOI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_5885_), .B(_5890_), .C(_5828_), .Y(_5891_) );
	OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_5529_), .B(_5891_), .C(_5820_), .Y(_5892_) );
	NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_5816_), .B(_5892_), .Y(_5893_) );
	NAND3X1 NAND3X1_1264 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf4), .B(_5845_), .C(_5893_), .Y(_5894_) );
	OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf3), .B(_5848_), .Y(_5895_) );
	NAND3X1 NAND3X1_1265 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf2), .B(_5895_), .C(_5894_), .Y(_5896_) );
	NAND3X1 NAND3X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_5815_), .B(_5896_), .C(_5889_), .Y(_5897_) );
	NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_5525_), .B(_5529_), .Y(_5898_) );
	INVX1 INVX1_946 ( .gnd(gnd), .vdd(vdd), .A(_5517_), .Y(_5900_) );
	AOI21X1 AOI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_5381_), .B(_5384_), .C(divider_absoluteValue_B_flipSign_result_22_bF_buf1), .Y(_5901_) );
	AOI21X1 AOI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_5901_), .B(_5523_), .C(_5900_), .Y(_5902_) );
	OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_5525_), .B(_5820_), .C(_5902_), .Y(_5903_) );
	AOI21X1 AOI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_5898_), .B(_5828_), .C(_5903_), .Y(_5904_) );
	AOI21X1 AOI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_5672_), .B(_5677_), .C(_5615_), .Y(_5905_) );
	OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_5838_), .B(_5905_), .C(_5545_), .Y(_5906_) );
	NAND3X1 NAND3X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_5904_), .B(_5906_), .C(_5813_), .Y(_5907_) );
	NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_5907_), .Y(_5908_) );
	OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .B(_5423_), .C(_5908_), .Y(_5909_) );
	NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_5419_), .B(_5424_), .Y(_5911_) );
	INVX1 INVX1_947 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .Y(_5912_) );
	OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_5828_), .B(_5841_), .C(_5528_), .Y(_5913_) );
	AOI21X1 AOI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(_5428_), .C(_5912_), .Y(_5914_) );
	NAND3X1 NAND3X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_5912_), .B(_5428_), .C(_5913_), .Y(_5915_) );
	INVX1 INVX1_948 ( .gnd(gnd), .vdd(vdd), .A(_5915_), .Y(_5916_) );
	OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_5914_), .B(_5916_), .C(divider_divuResult_8_bF_buf2), .Y(_5917_) );
	NAND3X1 NAND3X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf0), .B(_5909_), .C(_5917_), .Y(_5918_) );
	INVX1 INVX1_949 ( .gnd(gnd), .vdd(vdd), .A(_5909_), .Y(_5919_) );
	AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_5792_), .Y(_5920_) );
	OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_5693_), .B(_5920_), .C(_5890_), .Y(_5922_) );
	AOI21X1 AOI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_5922_), .B(_5511_), .C(_5434_), .Y(_5923_) );
	OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5923_), .C(_5911_), .Y(_5924_) );
	AOI21X1 AOI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_5924_), .B(_5915_), .C(_5908_), .Y(_5925_) );
	OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_5919_), .B(_5925_), .C(divider_absoluteValue_B_flipSign_result_22_bF_buf0), .Y(_5926_) );
	OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_5393_), .B(divider_divuResult_9_bF_buf3), .C(_5426_), .Y(_5927_) );
	NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_5434_), .B(_5891_), .Y(_5928_) );
	NAND3X1 NAND3X1_1270 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf1), .B(_5913_), .C(_5928_), .Y(_5929_) );
	OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_5927_), .B(divider_divuResult_8_bF_buf0), .C(_5929_), .Y(_5930_) );
	NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf3), .B(_5930_), .Y(_5931_) );
	OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf6), .B(_5927_), .Y(_5933_) );
	NAND3X1 NAND3X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf2), .B(_5929_), .C(_5933_), .Y(_5934_) );
	NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_5934_), .B(_5931_), .Y(_5935_) );
	NAND3X1 NAND3X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_5918_), .B(_5926_), .C(_5935_), .Y(_5936_) );
	NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_5897_), .B(_5936_), .Y(_5937_) );
	OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_5439_), .B(divider_divuResult_9_bF_buf2), .C(_5454_), .Y(_5938_) );
	OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf1), .B(_5886__bF_buf2), .C(_5938_), .Y(_5939_) );
	INVX1 INVX1_950 ( .gnd(gnd), .vdd(vdd), .A(_5543_), .Y(_5940_) );
	AOI21X1 AOI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_5840_), .B(_5839_), .C(_5940_), .Y(_5941_) );
	OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_5506_), .B(_5941_), .C(_5531_), .Y(_5942_) );
	NAND3X1 NAND3X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_5530_), .B(_5509_), .C(_5942_), .Y(_5944_) );
	INVX1 INVX1_951 ( .gnd(gnd), .vdd(vdd), .A(_5530_), .Y(_5945_) );
	OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_5693_), .B(_5920_), .C(_5543_), .Y(_5946_) );
	AOI22X1 AOI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_5467_), .B(_5469_), .C(_5824_), .D(_5946_), .Y(_5947_) );
	OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_5826_), .B(_5947_), .C(_5945_), .Y(_5948_) );
	NAND3X1 NAND3X1_1274 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf5), .B(_5944_), .C(_5948_), .Y(_5949_) );
	NAND3X1 NAND3X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf2), .B(_5939_), .C(_5949_), .Y(_5950_) );
	INVX1 INVX1_952 ( .gnd(gnd), .vdd(vdd), .A(_5938_), .Y(_5951_) );
	OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf0), .B(_5886__bF_buf1), .C(_5951_), .Y(_5952_) );
	OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_5826_), .B(_5947_), .C(_5530_), .Y(_5953_) );
	NAND3X1 NAND3X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_5945_), .B(_5509_), .C(_5942_), .Y(_5955_) );
	NAND3X1 NAND3X1_1277 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf4), .B(_5955_), .C(_5953_), .Y(_5956_) );
	NAND3X1 NAND3X1_1278 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf1), .B(_5952_), .C(_5956_), .Y(_5957_) );
	NOR3X1 NOR3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_5531_), .B(_5506_), .C(_5941_), .Y(_5958_) );
	OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_5958_), .B(_5947_), .C(divider_divuResult_8_bF_buf3), .Y(_5959_) );
	OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_5016_), .B(divider_divuResult_9_bF_buf1), .C(_5465_), .Y(_5960_) );
	OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf3), .B(_5886__bF_buf0), .C(_5960_), .Y(_5961_) );
	NAND3X1 NAND3X1_1279 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf0), .B(_5961_), .C(_5959_), .Y(_5962_) );
	INVX1 INVX1_953 ( .gnd(gnd), .vdd(vdd), .A(_5531_), .Y(_5963_) );
	NAND3X1 NAND3X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_5963_), .B(_5824_), .C(_5946_), .Y(_5964_) );
	AOI21X1 AOI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_5964_), .B(_5942_), .C(_5908_), .Y(_5965_) );
	INVX1 INVX1_954 ( .gnd(gnd), .vdd(vdd), .A(_5960_), .Y(_5966_) );
	NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_5966_), .B(divider_divuResult_8_bF_buf2), .Y(_5967_) );
	OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_5967_), .B(_5965_), .C(_3789__bF_buf4), .Y(_5968_) );
	NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_5962_), .B(_5968_), .Y(_5969_) );
	NAND3X1 NAND3X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_5969_), .B(_5950_), .C(_5957_), .Y(_5970_) );
	INVX1 INVX1_955 ( .gnd(gnd), .vdd(vdd), .A(_5535_), .Y(_5971_) );
	NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_5532_), .B(_5533_), .Y(_5972_) );
	INVX1 INVX1_956 ( .gnd(gnd), .vdd(vdd), .A(_5885_), .Y(_5973_) );
	NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_5542_), .B(_5973_), .Y(_5974_) );
	OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_5971_), .B(_5974_), .C(_5972_), .Y(_5977_) );
	INVX1 INVX1_957 ( .gnd(gnd), .vdd(vdd), .A(_5972_), .Y(_5978_) );
	OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_5973_), .B(_5542_), .Y(_5979_) );
	NAND3X1 NAND3X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_5535_), .B(_5978_), .C(_5979_), .Y(_5980_) );
	NAND3X1 NAND3X1_1283 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf1), .B(_5977_), .C(_5980_), .Y(_5981_) );
	OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_5473_), .B(divider_divuResult_9_bF_buf0), .C(_5489_), .Y(_5982_) );
	OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf0), .B(_5982_), .Y(_5983_) );
	AOI21X1 AOI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_5981_), .B(_5983_), .C(divider_absoluteValue_B_flipSign_result_18_bF_buf4), .Y(_5984_) );
	OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf6), .B(_5503_), .Y(_5985_) );
	XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_5885_), .B(_5542_), .Y(_5986_) );
	OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_5986_), .B(_5908_), .Y(_5988_) );
	AOI21X1 AOI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_5988_), .B(_5985_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf0), .Y(_5989_) );
	NAND3X1 NAND3X1_1284 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf3), .B(_5983_), .C(_5981_), .Y(_5990_) );
	AOI21X1 AOI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_5989_), .B(_5990_), .C(_5984_), .Y(_5991_) );
	AOI21X1 AOI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_5956_), .B(_5952_), .C(divider_absoluteValue_B_flipSign_result_20_bF_buf0), .Y(_5992_) );
	OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_5966_), .B(divider_divuResult_8_bF_buf5), .C(_5959_), .Y(_5993_) );
	NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf4), .B(_5993_), .Y(_5994_) );
	AOI21X1 AOI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_5957_), .B(_5994_), .C(_5992_), .Y(_5995_) );
	OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_5970_), .B(_5991_), .C(_5995_), .Y(_5996_) );
	NOR3X1 NOR3X1_57 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf3), .B(_5919_), .C(_5925_), .Y(_5997_) );
	NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf1), .B(_5930_), .Y(_5999_) );
	INVX1 INVX1_958 ( .gnd(gnd), .vdd(vdd), .A(_5999_), .Y(_6000_) );
	AOI21X1 AOI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_5926_), .B(_6000_), .C(_5997_), .Y(_6001_) );
	INVX1 INVX1_959 ( .gnd(gnd), .vdd(vdd), .A(_5814_), .Y(_6002_) );
	NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf0), .B(_6002_), .Y(_6003_) );
	AOI21X1 AOI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_5894_), .B(_5895_), .C(divider_absoluteValue_B_flipSign_result_23_bF_buf1), .Y(_6004_) );
	AOI21X1 AOI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_6004_), .B(_5815_), .C(_6003_), .Y(_6005_) );
	OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_5897_), .B(_6001_), .C(_6005_), .Y(_6006_) );
	AOI21X1 AOI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_5937_), .B(_5996_), .C(_6006_), .Y(_6007_) );
	AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_5950_), .B(_5957_), .Y(_6008_) );
	OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf2), .B(_5886__bF_buf3), .C(_5982_), .Y(_6010_) );
	OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_5971_), .B(_5974_), .C(_5978_), .Y(_6011_) );
	NAND3X1 NAND3X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_5535_), .B(_5972_), .C(_5979_), .Y(_6012_) );
	NAND3X1 NAND3X1_1286 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf4), .B(_6011_), .C(_6012_), .Y(_6013_) );
	NAND3X1 NAND3X1_1287 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf2), .B(_6010_), .C(_6013_), .Y(_6014_) );
	NAND3X1 NAND3X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf2), .B(_5983_), .C(_5981_), .Y(_6015_) );
	OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_5908_), .B(_5986_), .C(_5985_), .Y(_6016_) );
	NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .B(_6016_), .Y(_6017_) );
	NAND3X1 NAND3X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf4), .B(_5985_), .C(_5988_), .Y(_6018_) );
	AOI22X1 AOI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_6017_), .B(_6018_), .C(_6014_), .D(_6015_), .Y(_6019_) );
	NAND3X1 NAND3X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_5969_), .B(_6019_), .C(_6008_), .Y(_6020_) );
	NOR3X1 NOR3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_5897_), .B(_5936_), .C(_6020_), .Y(_6021_) );
	NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_5562_), .B(_5568_), .Y(_6022_) );
	INVX1 INVX1_960 ( .gnd(gnd), .vdd(vdd), .A(_5794_), .Y(_6023_) );
	OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .B(_5687_), .C(_5587_), .Y(_6024_) );
	OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_5810_), .B(_5882_), .C(_5678_), .Y(_6025_) );
	AOI22X1 AOI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_5836_), .B(_6024_), .C(_5613_), .D(_6025_), .Y(_6026_) );
	OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_6023_), .B(_6026_), .C(_5683_), .Y(_6027_) );
	NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_6022_), .B(_6027_), .Y(_6028_) );
	INVX1 INVX1_961 ( .gnd(gnd), .vdd(vdd), .A(_6022_), .Y(_6029_) );
	NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_5883_), .B(_5792_), .Y(_6032_) );
	AOI21X1 AOI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_6032_), .B(_5678_), .C(_5798_), .Y(_6033_) );
	OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_5690_), .B(_6033_), .C(_5794_), .Y(_6034_) );
	NAND3X1 NAND3X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_6029_), .B(_5683_), .C(_6034_), .Y(_6035_) );
	NAND3X1 NAND3X1_1292 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf3), .B(_6035_), .C(_6028_), .Y(_6036_) );
	OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_5563_), .B(divider_divuResult_9_bF_buf5), .C(_5561_), .Y(_6037_) );
	OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf2), .B(_6037_), .Y(_6038_) );
	AOI21X1 AOI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_6036_), .B(_6038_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf2), .Y(_6039_) );
	OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf1), .B(_5886__bF_buf2), .C(_6037_), .Y(_6040_) );
	NAND3X1 NAND3X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_6022_), .B(_5683_), .C(_6034_), .Y(_6041_) );
	OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_5831_), .B(_5681_), .C(_6027_), .Y(_6043_) );
	NAND3X1 NAND3X1_1294 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf1), .B(_6041_), .C(_6043_), .Y(_6044_) );
	AOI21X1 AOI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_6044_), .B(_6040_), .C(_2922__bF_buf0), .Y(_6045_) );
	NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_6023_), .B(_6026_), .Y(_6046_) );
	NOR3X1 NOR3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_5794_), .B(_5690_), .C(_6033_), .Y(_6047_) );
	OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_6047_), .B(_6046_), .C(divider_divuResult_8_bF_buf0), .Y(_6048_) );
	OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf0), .B(_5886__bF_buf1), .C(_5682_), .Y(_6049_) );
	NAND3X1 NAND3X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf4), .B(_6049_), .C(_6048_), .Y(_6050_) );
	NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_6023_), .B(_6026_), .Y(_6051_) );
	NAND3X1 NAND3X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_6034_), .B(_6051_), .C(divider_divuResult_8_bF_buf6), .Y(_6052_) );
	OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf5), .B(_5682_), .Y(_6054_) );
	NAND3X1 NAND3X1_1297 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .B(_6052_), .C(_6054_), .Y(_6055_) );
	NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_6050_), .B(_6055_), .Y(_6056_) );
	NOR3X1 NOR3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_6056_), .B(_6039_), .C(_6045_), .Y(_6057_) );
	NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_5796_), .B(_6025_), .Y(_6058_) );
	NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_6058_), .Y(_6059_) );
	NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_5797_), .B(_6059_), .Y(_6060_) );
	INVX1 INVX1_962 ( .gnd(gnd), .vdd(vdd), .A(_5797_), .Y(_6061_) );
	NAND3X1 NAND3X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_6061_), .C(_6058_), .Y(_6062_) );
	AOI21X1 AOI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_6060_), .B(_6062_), .C(_5908_), .Y(_6063_) );
	OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf3), .B(_5886__bF_buf0), .C(_5687_), .Y(_6065_) );
	INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_6065_), .Y(_6066_) );
	NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_6066_), .B(_6063_), .Y(_6067_) );
	NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf1), .B(_6067_), .Y(_6068_) );
	NAND3X1 NAND3X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_5797_), .C(_6058_), .Y(_6069_) );
	NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_6061_), .B(_6059_), .Y(_6070_) );
	NAND3X1 NAND3X1_1300 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf4), .B(_6069_), .C(_6070_), .Y(_6071_) );
	AOI21X1 AOI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_6071_), .B(_6065_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf0), .Y(_6072_) );
	INVX1 INVX1_963 ( .gnd(gnd), .vdd(vdd), .A(_6072_), .Y(_6073_) );
	XNOR2X1 XNOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .B(_5595_), .Y(_6074_) );
	AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf3), .B(_6074_), .Y(_6076_) );
	OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_5377__bF_buf3), .B(_5583_), .C(_5589_), .Y(_6077_) );
	INVX1 INVX1_964 ( .gnd(gnd), .vdd(vdd), .A(_6077_), .Y(_6078_) );
	NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_6078_), .B(divider_divuResult_8_bF_buf2), .Y(_6079_) );
	OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_6079_), .B(_6076_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .Y(_6080_) );
	NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_6074_), .B(divider_divuResult_8_bF_buf1), .Y(_6081_) );
	OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf2), .B(_5886__bF_buf3), .C(_6077_), .Y(_6082_) );
	NAND3X1 NAND3X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf3), .B(_6082_), .C(_6081_), .Y(_6083_) );
	AOI22X1 AOI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(_6080_), .B(_6083_), .C(_6073_), .D(_6068_), .Y(_6084_) );
	INVX1 INVX1_965 ( .gnd(gnd), .vdd(vdd), .A(_5646_), .Y(_6085_) );
	AOI21X1 AOI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_5792_), .B(_5809_), .C(_5671_), .Y(_6087_) );
	OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_6085_), .B(_6087_), .C(_5641_), .Y(_6088_) );
	NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .B(_6088_), .Y(_6089_) );
	INVX1 INVX1_966 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .Y(_6090_) );
	INVX1 INVX1_967 ( .gnd(gnd), .vdd(vdd), .A(_5809_), .Y(_6091_) );
	NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_6091_), .B(_5882_), .Y(_6092_) );
	OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_5671_), .B(_6092_), .C(_5648_), .Y(_6093_) );
	NAND3X1 NAND3X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_5641_), .B(_6090_), .C(_6093_), .Y(_6094_) );
	NAND3X1 NAND3X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_6089_), .B(_6094_), .C(divider_divuResult_8_bF_buf0), .Y(_6095_) );
	NAND3X1 NAND3X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_5616_), .B(_5626_), .C(_5908_), .Y(_6096_) );
	NAND3X1 NAND3X1_1305 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .B(_6096_), .C(_6095_), .Y(_6098_) );
	AOI21X1 AOI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_6095_), .B(_6096_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .Y(_6099_) );
	OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_5676_), .B(_6085_), .C(_6087_), .Y(_6100_) );
	NAND3X1 NAND3X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_6093_), .B(_6100_), .C(divider_divuResult_8_bF_buf6), .Y(_6101_) );
	NAND3X1 NAND3X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_5639_), .B(_5640_), .C(_5908_), .Y(_6102_) );
	AOI21X1 AOI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_6102_), .B(_6101_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .Y(_6103_) );
	OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_6103_), .B(_6099_), .C(_6098_), .Y(_6104_) );
	AOI21X1 AOI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_6095_), .B(_6096_), .C(_1484__bF_buf3), .Y(_6105_) );
	OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf1), .B(_5886__bF_buf2), .C(_5673_), .Y(_6106_) );
	NAND3X1 NAND3X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .B(_5641_), .C(_6093_), .Y(_6107_) );
	NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_6090_), .B(_6088_), .Y(_6109_) );
	NAND3X1 NAND3X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_6109_), .B(_6107_), .C(divider_divuResult_8_bF_buf5), .Y(_6110_) );
	AOI21X1 AOI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_6110_), .B(_6106_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .Y(_6111_) );
	AOI21X1 AOI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_6102_), .B(_6101_), .C(_1265__bF_buf0), .Y(_6112_) );
	NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_6100_), .B(_6093_), .Y(_6113_) );
	NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_6113_), .B(divider_divuResult_8_bF_buf4), .Y(_6114_) );
	NAND3X1 NAND3X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_5643_), .B(_5645_), .C(_5908_), .Y(_6115_) );
	AOI21X1 AOI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_6115_), .B(_6114_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .Y(_6116_) );
	OAI22X1 OAI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_6112_), .B(_6116_), .C(_6105_), .D(_6111_), .Y(_6117_) );
	OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_5800_), .B(_5802_), .C(_5908_), .Y(_6118_) );
	NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_5799_), .B(_5803_), .Y(_6120_) );
	NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_5804_), .B(_5808_), .Y(_6121_) );
	INVX1 INVX1_968 ( .gnd(gnd), .vdd(vdd), .A(_6121_), .Y(_6122_) );
	OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_6122_), .B(_5882_), .C(_5670_), .Y(_6123_) );
	NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_6120_), .B(_6123_), .Y(_6124_) );
	INVX1 INVX1_969 ( .gnd(gnd), .vdd(vdd), .A(_6120_), .Y(_6125_) );
	NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_6121_), .B(_5792_), .Y(_6126_) );
	NAND3X1 NAND3X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_5670_), .B(_6125_), .C(_6126_), .Y(_6127_) );
	NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_6127_), .B(_6124_), .Y(_6128_) );
	NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_6128_), .B(divider_divuResult_8_bF_buf3), .Y(_6129_) );
	NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_6129_), .B(_6118_), .Y(_6131_) );
	NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .B(_6131_), .Y(_6132_) );
	NAND3X1 NAND3X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_5662_), .B(_5663_), .C(_5908_), .Y(_6133_) );
	NAND3X1 NAND3X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_6124_), .B(_6127_), .C(divider_divuResult_8_bF_buf2), .Y(_6134_) );
	AOI21X1 AOI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_6133_), .B(_6134_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .Y(_6135_) );
	NAND3X1 NAND3X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_5667_), .B(_5668_), .C(_5908_), .Y(_6136_) );
	NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_6122_), .B(_5882_), .Y(_6137_) );
	NAND3X1 NAND3X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_6126_), .B(_6137_), .C(divider_divuResult_8_bF_buf1), .Y(_6138_) );
	AOI21X1 AOI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_6136_), .B(_6138_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .Y(_6139_) );
	OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .B(_6139_), .C(_6132_), .Y(_6140_) );
	OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_6140_), .B(_6117_), .C(_6104_), .Y(_6142_) );
	NAND3X1 NAND3X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_6084_), .B(_6142_), .C(_6057_), .Y(_6143_) );
	NAND3X1 NAND3X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf3), .B(_6040_), .C(_6044_), .Y(_6144_) );
	NAND3X1 NAND3X1_1318 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf1), .B(_6038_), .C(_6036_), .Y(_6145_) );
	NAND3X1 NAND3X1_1319 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .B(_6049_), .C(_6048_), .Y(_6146_) );
	NAND3X1 NAND3X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf3), .B(_6052_), .C(_6054_), .Y(_6147_) );
	NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_6146_), .B(_6147_), .Y(_6148_) );
	NAND3X1 NAND3X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_6145_), .B(_6144_), .C(_6148_), .Y(_6149_) );
	NOR3X1 NOR3X1_61 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .B(_6066_), .C(_6063_), .Y(_6150_) );
	OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_6066_), .B(_6063_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .Y(_6151_) );
	OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_6079_), .B(_6076_), .C(_1494__bF_buf2), .Y(_6153_) );
	INVX1 INVX1_970 ( .gnd(gnd), .vdd(vdd), .A(_6153_), .Y(_6154_) );
	AOI21X1 AOI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .B(_6151_), .C(_6150_), .Y(_6155_) );
	OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_6155_), .B(_6149_), .Y(_6156_) );
	INVX1 INVX1_971 ( .gnd(gnd), .vdd(vdd), .A(_6050_), .Y(_6157_) );
	AOI21X1 AOI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_6145_), .B(_6157_), .C(_6039_), .Y(_6158_) );
	NAND3X1 NAND3X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_6156_), .B(_6158_), .C(_6143_), .Y(_6159_) );
	NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_5859_), .B(divider_divuResult_8_bF_buf0), .Y(_6160_) );
	OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_5377__bF_buf2), .B(_5712_), .C(_5717_), .Y(_6161_) );
	INVX1 INVX1_972 ( .gnd(gnd), .vdd(vdd), .A(_6161_), .Y(_6162_) );
	INVX1 INVX1_973 ( .gnd(gnd), .vdd(vdd), .A(_5756_), .Y(_6164_) );
	OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_6164_), .B(_5791_), .C(_5858_), .Y(_6165_) );
	OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_5851_), .B(_5852_), .C(_6165_), .Y(_6166_) );
	OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_6162_), .C(_6166_), .Y(_6167_) );
	OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .B(_5850_), .C(_6167_), .Y(_6168_) );
	NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_5710_), .B(_5707_), .Y(_6169_) );
	OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_6167_), .B(_6169_), .Y(_6170_) );
	AOI21X1 AOI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_6168_), .B(_6170_), .C(_5908_), .Y(_6171_) );
	OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .B(_6171_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .Y(_6172_) );
	OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf0), .B(_5886__bF_buf1), .C(_5703_), .Y(_6173_) );
	AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_6167_), .B(_6169_), .Y(_6175_) );
	NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_6169_), .B(_6167_), .Y(_6176_) );
	OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_6175_), .B(_6176_), .C(divider_divuResult_8_bF_buf6), .Y(_6177_) );
	NAND3X1 NAND3X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_6173_), .C(_6177_), .Y(_6178_) );
	NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_5716_), .B(_5719_), .Y(_6179_) );
	XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_6165_), .B(_6179_), .Y(_6180_) );
	INVX1 INVX1_974 ( .gnd(gnd), .vdd(vdd), .A(_6180_), .Y(_6181_) );
	NAND3X1 NAND3X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6181_), .C(_5907_), .Y(_6182_) );
	OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf3), .B(_5886__bF_buf0), .C(_6162_), .Y(_6183_) );
	NAND3X1 NAND3X1_1325 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .B(_6182_), .C(_6183_), .Y(_6184_) );
	NAND3X1 NAND3X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6180_), .C(_5907_), .Y(_6186_) );
	OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf2), .B(_5886__bF_buf3), .C(_6161_), .Y(_6187_) );
	NAND3X1 NAND3X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf6), .B(_6186_), .C(_6187_), .Y(_6188_) );
	NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_6184_), .B(_6188_), .Y(_6189_) );
	NAND3X1 NAND3X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_6172_), .B(_6178_), .C(_6189_), .Y(_6190_) );
	NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_5747_), .B(_5751_), .Y(_6191_) );
	INVX1 INVX1_975 ( .gnd(gnd), .vdd(vdd), .A(_5752_), .Y(_6192_) );
	INVX1 INVX1_976 ( .gnd(gnd), .vdd(vdd), .A(_5755_), .Y(_6193_) );
	OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_6192_), .B(_6193_), .C(_5881_), .Y(_6194_) );
	AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_6194_), .B(_5741_), .Y(_6195_) );
	XNOR2X1 XNOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_6195_), .B(_6191_), .Y(_6197_) );
	OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf1), .B(_5886__bF_buf2), .C(_5854_), .Y(_6198_) );
	OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_5908_), .B(_6197_), .C(_6198_), .Y(_6199_) );
	NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .B(_6199_), .Y(_6200_) );
	OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf0), .B(_5886__bF_buf1), .C(_5856_), .Y(_6201_) );
	NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_6197_), .B(divider_divuResult_8_bF_buf5), .Y(_6202_) );
	AOI21X1 AOI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_6202_), .B(_6201_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .Y(_6203_) );
	OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_5739_), .B(divider_divuResult_9_bF_buf4), .C(_5754_), .Y(_6204_) );
	OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf3), .B(_5886__bF_buf0), .C(_6204_), .Y(_6205_) );
	NAND3X1 NAND3X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_5752_), .B(_5755_), .C(_5791_), .Y(_6206_) );
	NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_6206_), .B(_6194_), .Y(_6208_) );
	INVX1 INVX1_977 ( .gnd(gnd), .vdd(vdd), .A(_6208_), .Y(_6209_) );
	NAND3X1 NAND3X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6209_), .C(_5907_), .Y(_6210_) );
	AOI21X1 AOI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_6205_), .B(_6210_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .Y(_6211_) );
	OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_6211_), .B(_6203_), .C(_6200_), .Y(_6212_) );
	OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_5859_), .B(divider_divuResult_8_bF_buf4), .C(_6177_), .Y(_6213_) );
	INVX1 INVX1_978 ( .gnd(gnd), .vdd(vdd), .A(_6213_), .Y(_6214_) );
	OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_6161_), .B(divider_divuResult_8_bF_buf3), .C(_6182_), .Y(_6215_) );
	OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .B(_6215_), .C(_6178_), .Y(_6216_) );
	OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf2), .B(_6214_), .C(_6216_), .Y(_6217_) );
	OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_6212_), .B(_6190_), .C(_6217_), .Y(_6219_) );
	OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_5908_), .B(_6197_), .Y(_6220_) );
	NAND3X1 NAND3X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf2), .B(_6198_), .C(_6220_), .Y(_6221_) );
	NAND3X1 NAND3X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6208_), .C(_5907_), .Y(_6222_) );
	INVX1 INVX1_979 ( .gnd(gnd), .vdd(vdd), .A(_6204_), .Y(_6223_) );
	OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf2), .B(_5886__bF_buf3), .C(_6223_), .Y(_6224_) );
	NAND3X1 NAND3X1_1333 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(_6222_), .C(_6224_), .Y(_6225_) );
	NAND3X1 NAND3X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf1), .B(_6210_), .C(_6205_), .Y(_6226_) );
	NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_6225_), .B(_6226_), .Y(_6227_) );
	NAND3X1 NAND3X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_6200_), .B(_6221_), .C(_6227_), .Y(_6228_) );
	NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_6190_), .B(_6228_), .Y(_6230_) );
	OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf1), .B(_5886__bF_buf2), .C(_5864_), .Y(_6231_) );
	NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_5774_), .B(_5777_), .Y(_6232_) );
	NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_5871_), .B(_5872_), .Y(_6233_) );
	OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_6233_), .B(_5880_), .C(_5772_), .Y(_6234_) );
	XNOR2X1 XNOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_6234_), .B(_6232_), .Y(_6235_) );
	NAND3X1 NAND3X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6235_), .C(_5907_), .Y(_6236_) );
	NAND3X1 NAND3X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_6236_), .C(_6231_), .Y(_6237_) );
	INVX1 INVX1_980 ( .gnd(gnd), .vdd(vdd), .A(_6237_), .Y(_6238_) );
	INVX1 INVX1_981 ( .gnd(gnd), .vdd(vdd), .A(_5864_), .Y(_6239_) );
	OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_6239_), .B(divider_divuResult_8_bF_buf2), .C(_6236_), .Y(_6241_) );
	NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .B(_6241_), .Y(_6242_) );
	OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_5781_), .B(divider_divuResult_9_bF_buf3), .C(_5769_), .Y(_6243_) );
	INVX1 INVX1_982 ( .gnd(gnd), .vdd(vdd), .A(_6243_), .Y(_6244_) );
	OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf0), .B(_5886__bF_buf1), .C(_6244_), .Y(_6245_) );
	OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_5871_), .B(_5872_), .C(_5789_), .Y(_6246_) );
	NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_6233_), .B(_5880_), .Y(_6247_) );
	NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_6246_), .B(_6247_), .Y(_6248_) );
	INVX1 INVX1_983 ( .gnd(gnd), .vdd(vdd), .A(_6248_), .Y(_6249_) );
	NAND3X1 NAND3X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6249_), .C(_5907_), .Y(_6250_) );
	AOI21X1 AOI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_6245_), .B(_6250_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .Y(_6252_) );
	AOI21X1 AOI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_6242_), .B(_6252_), .C(_6238_), .Y(_6253_) );
	NAND3X1 NAND3X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6248_), .C(_5907_), .Y(_6254_) );
	OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf3), .B(_5886__bF_buf0), .C(_6243_), .Y(_6255_) );
	NAND3X1 NAND3X1_1340 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .B(_6254_), .C(_6255_), .Y(_6256_) );
	NAND3X1 NAND3X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_6250_), .C(_6245_), .Y(_6257_) );
	NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_6256_), .B(_6257_), .Y(_6258_) );
	NAND3X1 NAND3X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_6237_), .B(_6242_), .C(_6258_), .Y(_6259_) );
	OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_5293_), .B(_5377__bF_buf1), .C(_5875_), .Y(_6260_) );
	NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_5787_), .B(_5879_), .Y(_6261_) );
	XNOR2X1 XNOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_6261_), .B(_5874_), .Y(_6263_) );
	INVX1 INVX1_984 ( .gnd(gnd), .vdd(vdd), .A(_6263_), .Y(_6264_) );
	NAND3X1 NAND3X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6264_), .C(_5907_), .Y(_6265_) );
	OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_6260_), .B(divider_divuResult_8_bF_buf1), .C(_6265_), .Y(_6266_) );
	NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_6266_), .Y(_6267_) );
	OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf2), .B(_5886__bF_buf3), .C(divider_aOp_abs_8_), .Y(_6268_) );
	NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_5280_), .B(_5282_), .Y(_6269_) );
	INVX1 INVX1_985 ( .gnd(gnd), .vdd(vdd), .A(_6269_), .Y(_6270_) );
	NAND3X1 NAND3X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6270_), .C(_5907_), .Y(_6271_) );
	AOI21X1 AOI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_6268_), .B(_6271_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .Y(_6272_) );
	NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_6266_), .Y(_6274_) );
	AOI21X1 AOI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_6267_), .B(_6272_), .C(_6274_), .Y(_6275_) );
	OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_6275_), .B(_6259_), .C(_6253_), .Y(_6276_) );
	AOI21X1 AOI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_6276_), .B(_6230_), .C(_6219_), .Y(_6277_) );
	NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_7_), .B(_1746__bF_buf4), .Y(_6278_) );
	INVX1 INVX1_986 ( .gnd(gnd), .vdd(vdd), .A(_6278_), .Y(_6279_) );
	NAND3X1 NAND3X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6269_), .C(_5907_), .Y(_6280_) );
	OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf1), .B(_5886__bF_buf2), .C(_5279_), .Y(_6281_) );
	NAND3X1 NAND3X1_1346 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_6280_), .C(_6281_), .Y(_6282_) );
	NAND3X1 NAND3X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_6271_), .C(_6268_), .Y(_6283_) );
	NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_6282_), .B(_6283_), .Y(_6285_) );
	INVX1 INVX1_987 ( .gnd(gnd), .vdd(vdd), .A(_6260_), .Y(_6286_) );
	NAND3X1 NAND3X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_6263_), .C(_5907_), .Y(_6287_) );
	OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_6286_), .B(divider_divuResult_8_bF_buf0), .C(_6287_), .Y(_6288_) );
	NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_6288_), .Y(_6289_) );
	NAND3X1 NAND3X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_6267_), .B(_6289_), .C(_6285_), .Y(_6290_) );
	NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .B(_6290_), .Y(_6291_) );
	NAND3X1 NAND3X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_6279_), .B(_6230_), .C(_6291_), .Y(_6292_) );
	NAND3X1 NAND3X1_1351 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .B(_6106_), .C(_6110_), .Y(_6293_) );
	NAND3X1 NAND3X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf2), .B(_6096_), .C(_6095_), .Y(_6294_) );
	NAND3X1 NAND3X1_1353 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .B(_6114_), .C(_6115_), .Y(_6296_) );
	NAND3X1 NAND3X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_6101_), .C(_6102_), .Y(_6297_) );
	AOI22X1 AOI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(_6297_), .B(_6296_), .C(_6293_), .D(_6294_), .Y(_6298_) );
	NAND3X1 NAND3X1_1355 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .B(_6129_), .C(_6118_), .Y(_6299_) );
	NAND3X1 NAND3X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf2), .B(_6134_), .C(_6133_), .Y(_6300_) );
	OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_5649_), .B(divider_divuResult_9_bF_buf2), .C(_5667_), .Y(_6301_) );
	NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_6301_), .B(divider_divuResult_8_bF_buf6), .Y(_6302_) );
	NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_6126_), .B(_6137_), .Y(_6303_) );
	NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_6303_), .B(_5908_), .Y(_6304_) );
	OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_6302_), .B(_6304_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .Y(_6305_) );
	NAND3X1 NAND3X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf6), .B(_6138_), .C(_6136_), .Y(_6307_) );
	AOI22X1 AOI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_6300_), .B(_6299_), .C(_6307_), .D(_6305_), .Y(_6308_) );
	NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_6298_), .B(_6308_), .Y(_6309_) );
	INVX1 INVX1_988 ( .gnd(gnd), .vdd(vdd), .A(_6309_), .Y(_6310_) );
	NAND3X1 NAND3X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_6084_), .B(_6057_), .C(_6310_), .Y(_6311_) );
	AOI21X1 AOI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_6277_), .B(_6292_), .C(_6311_), .Y(_6312_) );
	OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .B(_6312_), .C(_6021_), .Y(_6313_) );
	AOI21X1 AOI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_6313_), .B(_6007_), .C(_4008__bF_buf4), .Y(divider_divuResult_7_) );
	NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_2031_), .Y(_6314_) );
	INVX8 INVX8_39 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .Y(_6315_) );
	INVX1 INVX1_989 ( .gnd(gnd), .vdd(vdd), .A(_5897_), .Y(_6317_) );
	INVX1 INVX1_990 ( .gnd(gnd), .vdd(vdd), .A(_5936_), .Y(_6318_) );
	NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_6317_), .B(_6318_), .Y(_6319_) );
	INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .Y(_6320_) );
	AOI21X1 AOI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_5917_), .B(_5909_), .C(_4881__bF_buf3), .Y(_6321_) );
	OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_5999_), .B(_6321_), .C(_5918_), .Y(_6322_) );
	INVX1 INVX1_991 ( .gnd(gnd), .vdd(vdd), .A(_6005_), .Y(_6323_) );
	AOI21X1 AOI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_6317_), .B(_6322_), .C(_6323_), .Y(_6324_) );
	OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_6320_), .B(_6319_), .C(_6324_), .Y(_6325_) );
	NOR3X1 NOR3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf2), .B(_6066_), .C(_6063_), .Y(_6326_) );
	NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_6083_), .B(_6080_), .Y(_6328_) );
	OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_6072_), .B(_6326_), .C(_6328_), .Y(_6329_) );
	NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_6329_), .B(_6149_), .Y(_6330_) );
	OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_6149_), .B(_6155_), .C(_6158_), .Y(_6331_) );
	AOI21X1 AOI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_6330_), .B(_6142_), .C(_6331_), .Y(_6332_) );
	INVX1 INVX1_992 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_7_), .Y(_6333_) );
	AOI22X1 AOI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_6333_), .C(_6282_), .D(_6283_), .Y(_6334_) );
	NAND3X1 NAND3X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf2), .B(_6280_), .C(_6281_), .Y(_6335_) );
	OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .B(_6266_), .C(_6335_), .Y(_6336_) );
	OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_6336_), .B(_6334_), .C(_6267_), .Y(_6337_) );
	OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .B(_6337_), .C(_6253_), .Y(_6339_) );
	AOI21X1 AOI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_6339_), .B(_6230_), .C(_6219_), .Y(_6340_) );
	OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_6311_), .B(_6340_), .C(_6332_), .Y(_6341_) );
	AOI21X1 AOI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_6341_), .B(_6021_), .C(_6325_), .Y(_6342_) );
	OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf3), .B(_6342__bF_buf4), .C(_5814_), .Y(_6343_) );
	INVX1 INVX1_993 ( .gnd(gnd), .vdd(vdd), .A(_6343_), .Y(_6344_) );
	NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf1), .B(_6315__bF_buf5), .Y(_6345_) );
	OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf1), .B(_6344_), .C(divider_absoluteValue_B_flipSign_result_25_), .Y(_6346_) );
	OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_6002_), .B(divider_divuResult_7_bF_buf6), .C(_2229__bF_buf4), .Y(_6347_) );
	OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_6347_), .B(divider_absoluteValue_B_flipSign_result_25_), .Y(_6348_) );
	OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_5848_), .B(divider_divuResult_8_bF_buf5), .C(_5894_), .Y(_6350_) );
	NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf0), .B(_6350_), .Y(_6351_) );
	NAND3X1 NAND3X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf0), .B(_5895_), .C(_5894_), .Y(_6352_) );
	NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_6352_), .B(_6351_), .Y(_6353_) );
	INVX1 INVX1_994 ( .gnd(gnd), .vdd(vdd), .A(_6353_), .Y(_6354_) );
	INVX1 INVX1_995 ( .gnd(gnd), .vdd(vdd), .A(_6219_), .Y(_6355_) );
	OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_6228_), .B(_6190_), .Y(_6356_) );
	INVX1 INVX1_996 ( .gnd(gnd), .vdd(vdd), .A(_6253_), .Y(_6357_) );
	NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_6237_), .B(_6242_), .Y(_6358_) );
	AOI21X1 AOI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_6256_), .B(_6257_), .C(_6358_), .Y(_6359_) );
	NAND3X1 NAND3X1_1361 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .B(_6271_), .C(_6268_), .Y(_6361_) );
	NAND3X1 NAND3X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_6279_), .B(_6335_), .C(_6361_), .Y(_6362_) );
	OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_5279_), .B(divider_divuResult_8_bF_buf4), .C(_6271_), .Y(_6363_) );
	AOI22X1 AOI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_6288_), .B(_2547__bF_buf4), .C(_1768__bF_buf1), .D(_6363_), .Y(_6364_) );
	AOI22X1 AOI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_6266_), .C(_6364_), .D(_6362_), .Y(_6365_) );
	AOI21X1 AOI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .B(_6365_), .C(_6357_), .Y(_6366_) );
	OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_6356_), .B(_6366_), .C(_6355_), .Y(_6367_) );
	NOR3X1 NOR3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_6329_), .B(_6149_), .C(_6309_), .Y(_6368_) );
	NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_6368_), .B(_6367_), .Y(_6369_) );
	AOI21X1 AOI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_6369_), .B(_6332_), .C(_6020_), .Y(_6370_) );
	OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .B(_6370_), .C(_6318_), .Y(_6372_) );
	AOI21X1 AOI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_6372_), .B(_6001_), .C(_6354_), .Y(_6373_) );
	AOI21X1 AOI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_5981_), .B(_5983_), .C(_3263__bF_buf1), .Y(_6374_) );
	AOI21X1 AOI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_6013_), .B(_6010_), .C(divider_absoluteValue_B_flipSign_result_18_bF_buf1), .Y(_6375_) );
	NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_6018_), .B(_6017_), .Y(_6376_) );
	OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_6374_), .B(_6375_), .C(_6376_), .Y(_6377_) );
	NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_5970_), .B(_6377_), .Y(_6378_) );
	OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .B(_6312_), .C(_6378_), .Y(_6379_) );
	AOI21X1 AOI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_6379_), .B(_6320_), .C(_5936_), .Y(_6380_) );
	NOR3X1 NOR3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_6353_), .B(_6322_), .C(_6380_), .Y(_6381_) );
	OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_6373_), .B(_6381_), .C(divider_divuResult_7_bF_buf5), .Y(_6383_) );
	OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf4), .B(_6350_), .Y(_6384_) );
	NAND3X1 NAND3X1_1363 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf3), .B(_6384_), .C(_6383_), .Y(_6385_) );
	OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_6322_), .B(_6380_), .C(_6353_), .Y(_6386_) );
	NAND3X1 NAND3X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_6354_), .B(_6001_), .C(_6372_), .Y(_6387_) );
	NAND3X1 NAND3X1_1365 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf3), .B(_6387_), .C(_6386_), .Y(_6388_) );
	OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf2), .B(_6342__bF_buf3), .C(_6350_), .Y(_6389_) );
	NAND3X1 NAND3X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf2), .B(_6389_), .C(_6388_), .Y(_6390_) );
	AOI22X1 AOI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_6346_), .B(_6348_), .C(_6390_), .D(_6385_), .Y(_6391_) );
	NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_5909_), .B(_5917_), .Y(_6392_) );
	OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf1), .B(_6342__bF_buf2), .C(_6392_), .Y(_6393_) );
	NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_6321_), .B(_5997_), .Y(_6394_) );
	OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .B(_6370_), .C(_5935_), .Y(_6395_) );
	NAND3X1 NAND3X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_6394_), .B(_5999_), .C(_6395_), .Y(_6396_) );
	INVX1 INVX1_997 ( .gnd(gnd), .vdd(vdd), .A(_6394_), .Y(_6397_) );
	AOI22X1 AOI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_5931_), .B(_5934_), .C(_6320_), .D(_6379_), .Y(_6398_) );
	OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_6000_), .B(_6398_), .C(_6397_), .Y(_6399_) );
	NAND3X1 NAND3X1_1368 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf2), .B(_6396_), .C(_6399_), .Y(_6400_) );
	NAND3X1 NAND3X1_1369 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf3), .B(_6393_), .C(_6400_), .Y(_6401_) );
	INVX1 INVX1_998 ( .gnd(gnd), .vdd(vdd), .A(_6393_), .Y(_6402_) );
	NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_6378_), .B(_5937_), .Y(_6404_) );
	OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_6404_), .B(_6332_), .C(_6007_), .Y(_6405_) );
	NAND3X1 NAND3X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_6378_), .B(_6368_), .C(_5937_), .Y(_6406_) );
	NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_6340_), .B(_6406_), .Y(_6407_) );
	OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_6407_), .B(_6405_), .C(_1615__bF_buf0), .Y(_6408_) );
	OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_6000_), .B(_6398_), .C(_6394_), .Y(_6409_) );
	NAND3X1 NAND3X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_6397_), .B(_5999_), .C(_6395_), .Y(_6410_) );
	AOI21X1 AOI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(_6410_), .C(_6408_), .Y(_6411_) );
	OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_6402_), .B(_6411_), .C(_5516__bF_buf3), .Y(_6412_) );
	NOR3X1 NOR3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_5935_), .B(_5996_), .C(_6370_), .Y(_6413_) );
	OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_6398_), .B(_6413_), .C(divider_divuResult_7_bF_buf1), .Y(_6415_) );
	INVX1 INVX1_999 ( .gnd(gnd), .vdd(vdd), .A(_5930_), .Y(_6416_) );
	OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf0), .B(_6342__bF_buf1), .C(_6416_), .Y(_6417_) );
	NAND3X1 NAND3X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf2), .B(_6417_), .C(_6415_), .Y(_6418_) );
	OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf5), .B(_6342__bF_buf0), .C(_5930_), .Y(_6419_) );
	INVX1 INVX1_1000 ( .gnd(gnd), .vdd(vdd), .A(_5935_), .Y(_6420_) );
	NAND3X1 NAND3X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_6420_), .B(_6320_), .C(_6379_), .Y(_6421_) );
	NAND3X1 NAND3X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_6421_), .B(_6395_), .C(divider_divuResult_7_bF_buf0), .Y(_6422_) );
	NAND3X1 NAND3X1_1375 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf2), .B(_6419_), .C(_6422_), .Y(_6423_) );
	NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_6423_), .B(_6418_), .Y(_6424_) );
	AOI21X1 AOI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_6412_), .B(_6401_), .C(_6424_), .Y(_6426_) );
	NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_6391_), .B(_6426_), .Y(_6427_) );
	OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_5951_), .B(divider_divuResult_8_bF_buf3), .C(_5949_), .Y(_6428_) );
	OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf4), .B(_6342__bF_buf4), .C(_6428_), .Y(_6429_) );
	INVX1 INVX1_1001 ( .gnd(gnd), .vdd(vdd), .A(_5994_), .Y(_6430_) );
	INVX1 INVX1_1002 ( .gnd(gnd), .vdd(vdd), .A(_5991_), .Y(_6431_) );
	AOI21X1 AOI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_6369_), .B(_6332_), .C(_6377_), .Y(_6432_) );
	OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_6431_), .B(_6432_), .C(_5969_), .Y(_6433_) );
	NAND3X1 NAND3X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .B(_6430_), .C(_6433_), .Y(_6434_) );
	INVX1 INVX1_1003 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .Y(_6435_) );
	OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .B(_6312_), .C(_6019_), .Y(_6437_) );
	AOI22X1 AOI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_5962_), .B(_5968_), .C(_5991_), .D(_6437_), .Y(_6438_) );
	OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_5994_), .B(_6438_), .C(_6435_), .Y(_6439_) );
	NAND3X1 NAND3X1_1377 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf6), .B(_6434_), .C(_6439_), .Y(_6440_) );
	NAND3X1 NAND3X1_1378 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf2), .B(_6429_), .C(_6440_), .Y(_6441_) );
	INVX1 INVX1_1004 ( .gnd(gnd), .vdd(vdd), .A(_6428_), .Y(_6442_) );
	OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf3), .B(_6342__bF_buf3), .C(_6442_), .Y(_6443_) );
	OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_5994_), .B(_6438_), .C(_6008_), .Y(_6444_) );
	NAND3X1 NAND3X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_6435_), .B(_6430_), .C(_6433_), .Y(_6445_) );
	NAND3X1 NAND3X1_1380 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf5), .B(_6445_), .C(_6444_), .Y(_6446_) );
	NAND3X1 NAND3X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf0), .B(_6443_), .C(_6446_), .Y(_6448_) );
	INVX1 INVX1_1005 ( .gnd(gnd), .vdd(vdd), .A(_5969_), .Y(_6449_) );
	NAND3X1 NAND3X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_6449_), .B(_5991_), .C(_6437_), .Y(_6450_) );
	INVX1 INVX1_1006 ( .gnd(gnd), .vdd(vdd), .A(_6450_), .Y(_6451_) );
	OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_6438_), .B(_6451_), .C(divider_divuResult_7_bF_buf4), .Y(_6452_) );
	OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf2), .B(_6342__bF_buf2), .C(_5993_), .Y(_6453_) );
	NAND3X1 NAND3X1_1383 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf3), .B(_6453_), .C(_6452_), .Y(_6454_) );
	AOI21X1 AOI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_6433_), .B(_6450_), .C(_6408_), .Y(_6455_) );
	INVX1 INVX1_1007 ( .gnd(gnd), .vdd(vdd), .A(_5993_), .Y(_6456_) );
	NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_6456_), .B(divider_divuResult_7_bF_buf3), .Y(_6457_) );
	OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_6457_), .B(_6455_), .C(_4011__bF_buf1), .Y(_6459_) );
	AOI22X1 AOI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(_6454_), .B(_6459_), .C(_6441_), .D(_6448_), .Y(_6460_) );
	NAND3X1 NAND3X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_5981_), .B(_5983_), .C(_6408_), .Y(_6461_) );
	NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_6015_), .Y(_6462_) );
	INVX1 INVX1_1008 ( .gnd(gnd), .vdd(vdd), .A(_6462_), .Y(_6463_) );
	INVX1 INVX1_1009 ( .gnd(gnd), .vdd(vdd), .A(_6016_), .Y(_6464_) );
	OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .B(_6312_), .C(_6376_), .Y(_6465_) );
	OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .B(_6464_), .C(_6465_), .Y(_6466_) );
	NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_6463_), .B(_6466_), .Y(_6467_) );
	INVX1 INVX1_1010 ( .gnd(gnd), .vdd(vdd), .A(_5989_), .Y(_6468_) );
	NAND3X1 NAND3X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .B(_6462_), .C(_6465_), .Y(_6470_) );
	NAND3X1 NAND3X1_1386 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf2), .B(_6470_), .C(_6467_), .Y(_6471_) );
	NAND3X1 NAND3X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf3), .B(_6461_), .C(_6471_), .Y(_6472_) );
	AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_6341_), .B(_6376_), .Y(_6473_) );
	NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_6376_), .B(_6341_), .Y(_6474_) );
	OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_6473_), .B(_6474_), .C(divider_divuResult_7_bF_buf1), .Y(_6475_) );
	OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf1), .B(_6342__bF_buf1), .C(_6464_), .Y(_6476_) );
	NAND3X1 NAND3X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf0), .B(_6476_), .C(_6475_), .Y(_6477_) );
	AOI21X1 AOI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_6471_), .B(_6461_), .C(_3789__bF_buf2), .Y(_6478_) );
	OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .B(_6478_), .C(_6472_), .Y(_6479_) );
	NAND3X1 NAND3X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf3), .B(_6429_), .C(_6440_), .Y(_6481_) );
	AOI21X1 AOI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_6440_), .B(_6429_), .C(_4424__bF_buf2), .Y(_6482_) );
	NAND3X1 NAND3X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf0), .B(_6453_), .C(_6452_), .Y(_6483_) );
	OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .B(_6482_), .C(_6481_), .Y(_6484_) );
	AOI21X1 AOI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_6460_), .B(_6479_), .C(_6484_), .Y(_6485_) );
	NAND3X1 NAND3X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf2), .B(_6393_), .C(_6400_), .Y(_6486_) );
	AOI21X1 AOI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_6400_), .B(_6393_), .C(_5516__bF_buf1), .Y(_6487_) );
	OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .B(_6487_), .C(_6486_), .Y(_6488_) );
	AOI21X1 AOI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_6343_), .B(_2229__bF_buf3), .C(divider_absoluteValue_B_flipSign_result_25_), .Y(_6489_) );
	INVX1 INVX1_1011 ( .gnd(gnd), .vdd(vdd), .A(_6489_), .Y(_6490_) );
	NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_6347_), .Y(_6492_) );
	NAND3X1 NAND3X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf1), .B(_6384_), .C(_6383_), .Y(_6493_) );
	OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_6492_), .B(_6493_), .C(_6490_), .Y(_6494_) );
	AOI21X1 AOI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_6391_), .B(_6488_), .C(_6494_), .Y(_6495_) );
	OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_6427_), .B(_6485_), .C(_6495_), .Y(_6496_) );
	NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_6489_), .B(_6492_), .Y(_6497_) );
	NAND3X1 NAND3X1_1393 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf2), .B(_6389_), .C(_6388_), .Y(_6498_) );
	NAND3X1 NAND3X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_6497_), .B(_6498_), .C(_6493_), .Y(_6499_) );
	OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_6402_), .B(_6411_), .C(divider_absoluteValue_B_flipSign_result_23_bF_buf2), .Y(_6500_) );
	AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .B(_6423_), .Y(_6501_) );
	NAND3X1 NAND3X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_6486_), .B(_6500_), .C(_6501_), .Y(_6503_) );
	NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_6499_), .B(_6503_), .Y(_6504_) );
	NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_6441_), .B(_6448_), .Y(_6505_) );
	NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_6459_), .B(_6454_), .Y(_6506_) );
	NAND3X1 NAND3X1_1396 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf3), .B(_6461_), .C(_6471_), .Y(_6507_) );
	OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_6374_), .B(_6375_), .C(_6466_), .Y(_6508_) );
	NAND3X1 NAND3X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .B(_6463_), .C(_6465_), .Y(_6509_) );
	NAND3X1 NAND3X1_1398 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf0), .B(_6509_), .C(_6508_), .Y(_6510_) );
	OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(divider_divuResult_8_bF_buf2), .C(_5981_), .Y(_6511_) );
	OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf0), .B(_6342__bF_buf0), .C(_6511_), .Y(_6512_) );
	NAND3X1 NAND3X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf1), .B(_6512_), .C(_6510_), .Y(_6514_) );
	OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_6341_), .B(_6376_), .Y(_6515_) );
	NAND3X1 NAND3X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_6465_), .B(_6515_), .C(divider_divuResult_7_bF_buf6), .Y(_6516_) );
	OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf5), .B(_6342__bF_buf4), .C(_6016_), .Y(_6517_) );
	NAND3X1 NAND3X1_1401 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf0), .B(_6517_), .C(_6516_), .Y(_6518_) );
	NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .B(_6518_), .Y(_6519_) );
	AOI21X1 AOI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_6507_), .B(_6514_), .C(_6519_), .Y(_6520_) );
	NAND3X1 NAND3X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_6506_), .B(_6520_), .C(_6505_), .Y(_6521_) );
	INVX1 INVX1_1012 ( .gnd(gnd), .vdd(vdd), .A(_6521_), .Y(_6522_) );
	NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_6522_), .B(_6504_), .Y(_6523_) );
	NAND3X1 NAND3X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_6036_), .B(_6038_), .C(_6408_), .Y(_6525_) );
	NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_6039_), .B(_6045_), .Y(_6526_) );
	AOI21X1 AOI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .B(_6310_), .C(_6142_), .Y(_6527_) );
	OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_6329_), .B(_6527_), .C(_6155_), .Y(_6528_) );
	NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_6148_), .B(_6528_), .Y(_6529_) );
	NAND3X1 NAND3X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_6526_), .B(_6050_), .C(_6529_), .Y(_6530_) );
	INVX1 INVX1_1013 ( .gnd(gnd), .vdd(vdd), .A(_6526_), .Y(_6531_) );
	AOI21X1 AOI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_6277_), .B(_6292_), .C(_6309_), .Y(_6532_) );
	OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_6142_), .B(_6532_), .C(_6084_), .Y(_6533_) );
	AOI22X1 AOI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(_6146_), .B(_6147_), .C(_6155_), .D(_6533_), .Y(_6534_) );
	OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_6157_), .B(_6534_), .C(_6531_), .Y(_6536_) );
	NAND3X1 NAND3X1_1405 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf5), .B(_6530_), .C(_6536_), .Y(_6537_) );
	NAND3X1 NAND3X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf3), .B(_6525_), .C(_6537_), .Y(_6538_) );
	OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_6037_), .B(divider_divuResult_8_bF_buf1), .C(_6036_), .Y(_6539_) );
	OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf4), .B(_6342__bF_buf3), .C(_6539_), .Y(_6540_) );
	OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_6157_), .B(_6534_), .C(_6526_), .Y(_6541_) );
	NAND3X1 NAND3X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_6531_), .B(_6050_), .C(_6529_), .Y(_6542_) );
	NAND3X1 NAND3X1_1408 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf4), .B(_6542_), .C(_6541_), .Y(_6543_) );
	NAND3X1 NAND3X1_1409 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .B(_6540_), .C(_6543_), .Y(_6544_) );
	NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_6148_), .B(_6528_), .Y(_6545_) );
	OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_6534_), .B(_6545_), .C(divider_divuResult_7_bF_buf3), .Y(_6547_) );
	NAND3X1 NAND3X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_6052_), .B(_6054_), .C(_6408_), .Y(_6548_) );
	NAND3X1 NAND3X1_1411 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf0), .B(_6548_), .C(_6547_), .Y(_6549_) );
	NAND3X1 NAND3X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_6056_), .B(_6155_), .C(_6533_), .Y(_6550_) );
	NAND3X1 NAND3X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_6550_), .B(_6529_), .C(divider_divuResult_7_bF_buf2), .Y(_6551_) );
	OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_5682_), .B(divider_divuResult_8_bF_buf0), .C(_6052_), .Y(_6552_) );
	OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf3), .B(_6342__bF_buf2), .C(_6552_), .Y(_6553_) );
	NAND3X1 NAND3X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf2), .B(_6553_), .C(_6551_), .Y(_6554_) );
	NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_6554_), .B(_6549_), .Y(_6555_) );
	NAND3X1 NAND3X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_6538_), .B(_6544_), .C(_6555_), .Y(_6556_) );
	NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_6073_), .B(_6068_), .Y(_6558_) );
	OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_6142_), .B(_6532_), .C(_6328_), .Y(_6559_) );
	NAND3X1 NAND3X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .B(_6153_), .C(_6559_), .Y(_6560_) );
	INVX1 INVX1_1014 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .Y(_6561_) );
	INVX1 INVX1_1015 ( .gnd(gnd), .vdd(vdd), .A(_6328_), .Y(_6562_) );
	OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_6562_), .B(_6527_), .C(_6153_), .Y(_6563_) );
	OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_6150_), .B(_6561_), .C(_6563_), .Y(_6564_) );
	NAND3X1 NAND3X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(divider_divuResult_7_bF_buf1), .C(_6564_), .Y(_6565_) );
	OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_6063_), .B(_6066_), .C(_6408_), .Y(_6566_) );
	NAND3X1 NAND3X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf2), .B(_6566_), .C(_6565_), .Y(_6567_) );
	OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .B(_6072_), .C(_6563_), .Y(_6569_) );
	INVX1 INVX1_1016 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .Y(_6570_) );
	NAND3X1 NAND3X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_6570_), .B(_6153_), .C(_6559_), .Y(_6571_) );
	AOI21X1 AOI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_6569_), .B(_6571_), .C(_6408_), .Y(_6572_) );
	INVX1 INVX1_1017 ( .gnd(gnd), .vdd(vdd), .A(_6566_), .Y(_6573_) );
	OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_6572_), .B(_6573_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .Y(_6574_) );
	NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_6562_), .B(_6527_), .Y(_6575_) );
	NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_6559_), .B(_6575_), .Y(_6576_) );
	NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_6576_), .B(divider_divuResult_7_bF_buf0), .Y(_6577_) );
	NAND3X1 NAND3X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_6081_), .B(_6082_), .C(_6408_), .Y(_6578_) );
	NAND3X1 NAND3X1_1421 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .B(_6578_), .C(_6577_), .Y(_6580_) );
	NAND3X1 NAND3X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_6559_), .B(_6575_), .C(divider_divuResult_7_bF_buf6), .Y(_6581_) );
	OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_6078_), .B(divider_divuResult_8_bF_buf6), .C(_6081_), .Y(_6582_) );
	OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf2), .B(_6342__bF_buf1), .C(_6582_), .Y(_6583_) );
	NAND3X1 NAND3X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf1), .B(_6583_), .C(_6581_), .Y(_6584_) );
	NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_6580_), .B(_6584_), .Y(_6585_) );
	NAND3X1 NAND3X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_6567_), .B(_6574_), .C(_6585_), .Y(_6586_) );
	NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .B(_6556_), .Y(_6587_) );
	NAND3X1 NAND3X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_6095_), .B(_6096_), .C(_6408_), .Y(_6588_) );
	INVX1 INVX1_1018 ( .gnd(gnd), .vdd(vdd), .A(_6103_), .Y(_6589_) );
	NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .B(_6294_), .Y(_6591_) );
	NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_6296_), .B(_6297_), .Y(_6592_) );
	INVX1 INVX1_1019 ( .gnd(gnd), .vdd(vdd), .A(_6140_), .Y(_6593_) );
	INVX1 INVX1_1020 ( .gnd(gnd), .vdd(vdd), .A(_6308_), .Y(_6594_) );
	AOI21X1 AOI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_6277_), .B(_6292_), .C(_6594_), .Y(_6595_) );
	OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_6593_), .B(_6595_), .C(_6592_), .Y(_6596_) );
	NAND3X1 NAND3X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_6589_), .B(_6591_), .C(_6596_), .Y(_6597_) );
	INVX1 INVX1_1021 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6598_) );
	INVX1 INVX1_1022 ( .gnd(gnd), .vdd(vdd), .A(_6592_), .Y(_6599_) );
	AOI21X1 AOI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .B(_6308_), .C(_6593_), .Y(_6600_) );
	OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_6599_), .B(_6600_), .C(_6589_), .Y(_6602_) );
	NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_6598_), .B(_6602_), .Y(_6603_) );
	NAND3X1 NAND3X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_6597_), .B(_6603_), .C(divider_divuResult_7_bF_buf5), .Y(_6604_) );
	NAND3X1 NAND3X1_1428 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_6588_), .C(_6604_), .Y(_6605_) );
	OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_5673_), .B(divider_divuResult_8_bF_buf5), .C(_6095_), .Y(_6606_) );
	OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf1), .B(_6342__bF_buf0), .C(_6606_), .Y(_6607_) );
	OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_6105_), .B(_6111_), .C(_6602_), .Y(_6608_) );
	NAND3X1 NAND3X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_6589_), .B(_6598_), .C(_6596_), .Y(_6609_) );
	NAND3X1 NAND3X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_6609_), .B(divider_divuResult_7_bF_buf4), .C(_6608_), .Y(_6610_) );
	NAND3X1 NAND3X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf1), .B(_6607_), .C(_6610_), .Y(_6611_) );
	NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_6599_), .B(_6600_), .Y(_6613_) );
	NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_6596_), .B(_6613_), .Y(_6614_) );
	NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_6614_), .B(divider_divuResult_7_bF_buf3), .Y(_6615_) );
	NAND3X1 NAND3X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_6101_), .B(_6102_), .C(_6408_), .Y(_6616_) );
	NAND3X1 NAND3X1_1433 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .B(_6616_), .C(_6615_), .Y(_6617_) );
	AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_6613_), .B(_6596_), .Y(_6618_) );
	NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_6618_), .B(divider_divuResult_7_bF_buf2), .Y(_6619_) );
	NAND3X1 NAND3X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_6114_), .B(_6115_), .C(_6408_), .Y(_6620_) );
	NAND3X1 NAND3X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf1), .B(_6620_), .C(_6619_), .Y(_6621_) );
	AOI22X1 AOI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(_6617_), .B(_6621_), .C(_6605_), .D(_6611_), .Y(_6622_) );
	OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf0), .B(_6342__bF_buf4), .C(_6131_), .Y(_6624_) );
	NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_6021_), .B(_6159_), .Y(_6625_) );
	NAND3X1 NAND3X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .B(_6368_), .C(_6021_), .Y(_6626_) );
	NAND3X1 NAND3X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_6007_), .B(_6625_), .C(_6626_), .Y(_6627_) );
	INVX1 INVX1_1023 ( .gnd(gnd), .vdd(vdd), .A(_6135_), .Y(_6628_) );
	NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_6132_), .B(_6628_), .Y(_6629_) );
	INVX1 INVX1_1024 ( .gnd(gnd), .vdd(vdd), .A(_6629_), .Y(_6630_) );
	AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_6305_), .B(_6307_), .Y(_6631_) );
	AOI21X1 AOI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_6277_), .B(_6292_), .C(_6631_), .Y(_6632_) );
	OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_6139_), .B(_6632_), .C(_6630_), .Y(_6633_) );
	INVX1 INVX1_1025 ( .gnd(gnd), .vdd(vdd), .A(_6139_), .Y(_6635_) );
	INVX1 INVX1_1026 ( .gnd(gnd), .vdd(vdd), .A(_6631_), .Y(_6636_) );
	NAND2X1 NAND2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_6636_), .B(_6367_), .Y(_6637_) );
	NAND3X1 NAND3X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_6635_), .B(_6629_), .C(_6637_), .Y(_6638_) );
	NAND2X1 NAND2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_6638_), .B(_6633_), .Y(_6639_) );
	NAND3X1 NAND3X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf4), .B(_6627__bF_buf3), .C(_6639_), .Y(_6640_) );
	NAND3X1 NAND3X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf4), .B(_6624_), .C(_6640_), .Y(_6641_) );
	NAND2X1 NAND2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_6631_), .B(_6340_), .Y(_6642_) );
	NAND2X1 NAND2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_6637_), .B(_6642_), .Y(_6643_) );
	NAND3X1 NAND3X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf3), .B(_6643_), .C(_6627__bF_buf2), .Y(_6644_) );
	OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_6301_), .B(divider_divuResult_8_bF_buf4), .C(_6138_), .Y(_6646_) );
	INVX1 INVX1_1027 ( .gnd(gnd), .vdd(vdd), .A(_6646_), .Y(_6647_) );
	OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf5), .B(_6342__bF_buf3), .C(_6647_), .Y(_6648_) );
	NAND3X1 NAND3X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf1), .B(_6644_), .C(_6648_), .Y(_6649_) );
	AOI21X1 AOI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_6640_), .B(_6624_), .C(_1265__bF_buf3), .Y(_6650_) );
	OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_6650_), .C(_6641_), .Y(_6651_) );
	NAND3X1 NAND3X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf0), .B(_6588_), .C(_6604_), .Y(_6652_) );
	AOI21X1 AOI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_6604_), .B(_6588_), .C(_1494__bF_buf4), .Y(_6653_) );
	NAND3X1 NAND3X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf0), .B(_6616_), .C(_6615_), .Y(_6654_) );
	OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_6654_), .B(_6653_), .C(_6652_), .Y(_6655_) );
	AOI21X1 AOI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_6622_), .B(_6651_), .C(_6655_), .Y(_6657_) );
	INVX1 INVX1_1028 ( .gnd(gnd), .vdd(vdd), .A(_6657_), .Y(_6658_) );
	OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_6067_), .B(divider_divuResult_7_bF_buf1), .C(_6565_), .Y(_6659_) );
	INVX1 INVX1_1029 ( .gnd(gnd), .vdd(vdd), .A(_6659_), .Y(_6660_) );
	OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_6582_), .B(divider_divuResult_7_bF_buf0), .C(_6577_), .Y(_6661_) );
	OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf2), .B(_6661_), .C(_6567_), .Y(_6662_) );
	OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf1), .B(_6660_), .C(_6662_), .Y(_6663_) );
	AOI21X1 AOI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_6543_), .B(_6540_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .Y(_6664_) );
	NAND3X1 NAND3X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf1), .B(_6548_), .C(_6547_), .Y(_6665_) );
	INVX1 INVX1_1030 ( .gnd(gnd), .vdd(vdd), .A(_6665_), .Y(_6666_) );
	AOI21X1 AOI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(_6544_), .C(_6664_), .Y(_6668_) );
	OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_6663_), .B(_6556_), .C(_6668_), .Y(_6669_) );
	AOI21X1 AOI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_6587_), .B(_6658_), .C(_6669_), .Y(_6670_) );
	OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf4), .B(_6342__bF_buf2), .C(_6213_), .Y(_6671_) );
	AOI21X1 AOI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_6177_), .B(_6173_), .C(_7204__bF_buf1), .Y(_6672_) );
	INVX1 INVX1_1031 ( .gnd(gnd), .vdd(vdd), .A(_6178_), .Y(_6673_) );
	NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_6672_), .B(_6673_), .Y(_6674_) );
	NAND3X1 NAND3X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf5), .B(_6182_), .C(_6183_), .Y(_6675_) );
	NAND3X1 NAND3X1_1447 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_6186_), .C(_6187_), .Y(_6676_) );
	NAND2X1 NAND2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_6675_), .B(_6676_), .Y(_6677_) );
	INVX1 INVX1_1032 ( .gnd(gnd), .vdd(vdd), .A(_6212_), .Y(_6679_) );
	INVX1 INVX1_1033 ( .gnd(gnd), .vdd(vdd), .A(_6228_), .Y(_6680_) );
	AOI21X1 AOI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_6339_), .B(_6680_), .C(_6679_), .Y(_6681_) );
	OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_6677_), .B(_6681_), .C(_6675_), .Y(_6682_) );
	AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_6682_), .B(_6674_), .Y(_6683_) );
	NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_6674_), .B(_6682_), .Y(_6684_) );
	OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_6683_), .B(_6684_), .C(divider_divuResult_7_bF_buf6), .Y(_6685_) );
	NAND3X1 NAND3X1_1448 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_6671_), .C(_6685_), .Y(_6686_) );
	AOI21X1 AOI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_6627__bF_buf1), .B(_1615__bF_buf2), .C(_6214_), .Y(_6687_) );
	NAND2X1 NAND2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_6674_), .B(_6682_), .Y(_6688_) );
	OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_6682_), .B(_6674_), .Y(_6690_) );
	AOI21X1 AOI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_6688_), .B(_6690_), .C(_6408_), .Y(_6691_) );
	OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_6687_), .B(_6691_), .C(_8971__bF_buf5), .Y(_6692_) );
	NAND2X1 NAND2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_6686_), .B(_6692_), .Y(_6693_) );
	OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_6228_), .B(_6366_), .C(_6212_), .Y(_6694_) );
	NAND2X1 NAND2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_6189_), .B(_6694_), .Y(_6695_) );
	NAND2X1 NAND2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_6677_), .B(_6681_), .Y(_6696_) );
	NAND2X1 NAND2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_6695_), .B(_6696_), .Y(_6697_) );
	NAND3X1 NAND3X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf1), .B(_6697_), .C(_6627__bF_buf0), .Y(_6698_) );
	OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf3), .B(_6342__bF_buf1), .C(_6215_), .Y(_6699_) );
	NAND3X1 NAND3X1_1450 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .B(_6698_), .C(_6699_), .Y(_6701_) );
	INVX1 INVX1_1034 ( .gnd(gnd), .vdd(vdd), .A(_6697_), .Y(_6702_) );
	NAND3X1 NAND3X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf0), .B(_6702_), .C(_6627__bF_buf3), .Y(_6703_) );
	INVX1 INVX1_1035 ( .gnd(gnd), .vdd(vdd), .A(_6215_), .Y(_6704_) );
	OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf2), .B(_6342__bF_buf0), .C(_6704_), .Y(_6705_) );
	NAND3X1 NAND3X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf0), .B(_6703_), .C(_6705_), .Y(_6706_) );
	NAND2X1 NAND2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_6701_), .B(_6706_), .Y(_6707_) );
	OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf1), .B(_6342__bF_buf4), .C(_6199_), .Y(_6708_) );
	NAND2X1 NAND2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_6200_), .B(_6221_), .Y(_6709_) );
	INVX1 INVX1_1036 ( .gnd(gnd), .vdd(vdd), .A(_6211_), .Y(_6710_) );
	INVX1 INVX1_1037 ( .gnd(gnd), .vdd(vdd), .A(_6227_), .Y(_6712_) );
	OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_6712_), .B(_6366_), .C(_6710_), .Y(_6713_) );
	XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_6713_), .B(_6709_), .Y(_6714_) );
	NAND3X1 NAND3X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf4), .B(_6714_), .C(_6627__bF_buf2), .Y(_6715_) );
	NAND3X1 NAND3X1_1454 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(_6715_), .C(_6708_), .Y(_6716_) );
	INVX1 INVX1_1038 ( .gnd(gnd), .vdd(vdd), .A(_6199_), .Y(_6717_) );
	OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf0), .B(_6342__bF_buf3), .C(_6717_), .Y(_6718_) );
	XNOR2X1 XNOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_6713_), .B(_6709_), .Y(_6719_) );
	NAND3X1 NAND3X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf3), .B(_6719_), .C(_6627__bF_buf1), .Y(_6720_) );
	NAND3X1 NAND3X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf4), .B(_6720_), .C(_6718_), .Y(_6721_) );
	XNOR2X1 XNOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_6366_), .B(_6227_), .Y(_6723_) );
	INVX1 INVX1_1039 ( .gnd(gnd), .vdd(vdd), .A(_6723_), .Y(_6724_) );
	NAND3X1 NAND3X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf2), .B(_6724_), .C(_6627__bF_buf0), .Y(_6725_) );
	OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_6223_), .B(divider_divuResult_8_bF_buf3), .C(_6210_), .Y(_6726_) );
	INVX1 INVX1_1040 ( .gnd(gnd), .vdd(vdd), .A(_6726_), .Y(_6727_) );
	OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf5), .B(_6342__bF_buf2), .C(_6727_), .Y(_6728_) );
	NAND3X1 NAND3X1_1458 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .B(_6725_), .C(_6728_), .Y(_6729_) );
	OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf4), .B(_6342__bF_buf1), .C(_6726_), .Y(_6730_) );
	NAND3X1 NAND3X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf1), .B(_6723_), .C(_6627__bF_buf3), .Y(_6731_) );
	NAND3X1 NAND3X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_6731_), .C(_6730_), .Y(_6732_) );
	AOI22X1 AOI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(_6716_), .B(_6721_), .C(_6729_), .D(_6732_), .Y(_6734_) );
	NAND3X1 NAND3X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_6707_), .B(_6734_), .C(_6693_), .Y(_6735_) );
	OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf3), .B(_6342__bF_buf0), .C(_6241_), .Y(_6736_) );
	INVX1 INVX1_1041 ( .gnd(gnd), .vdd(vdd), .A(_6252_), .Y(_6737_) );
	INVX1 INVX1_1042 ( .gnd(gnd), .vdd(vdd), .A(_6258_), .Y(_6738_) );
	OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_6738_), .B(_6337_), .C(_6737_), .Y(_6739_) );
	XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_6739_), .B(_6358_), .Y(_6740_) );
	NAND3X1 NAND3X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf0), .B(_6740_), .C(_6627__bF_buf2), .Y(_6741_) );
	NAND3X1 NAND3X1_1463 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .B(_6741_), .C(_6736_), .Y(_6742_) );
	INVX1 INVX1_1043 ( .gnd(gnd), .vdd(vdd), .A(_6740_), .Y(_6743_) );
	NAND3X1 NAND3X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf4), .B(_6743_), .C(_6627__bF_buf1), .Y(_6745_) );
	INVX1 INVX1_1044 ( .gnd(gnd), .vdd(vdd), .A(_6241_), .Y(_6746_) );
	OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf2), .B(_6342__bF_buf4), .C(_6746_), .Y(_6747_) );
	NAND3X1 NAND3X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf0), .B(_6745_), .C(_6747_), .Y(_6748_) );
	XNOR2X1 XNOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_6365_), .B(_6738_), .Y(_6749_) );
	INVX1 INVX1_1045 ( .gnd(gnd), .vdd(vdd), .A(_6749_), .Y(_6750_) );
	NAND3X1 NAND3X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf3), .B(_6750_), .C(_6627__bF_buf0), .Y(_6751_) );
	OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_6243_), .B(divider_divuResult_8_bF_buf2), .C(_6250_), .Y(_6752_) );
	INVX1 INVX1_1046 ( .gnd(gnd), .vdd(vdd), .A(_6752_), .Y(_6753_) );
	OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf1), .B(_6342__bF_buf3), .C(_6753_), .Y(_6754_) );
	NAND3X1 NAND3X1_1467 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .B(_6751_), .C(_6754_), .Y(_6756_) );
	NAND3X1 NAND3X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf2), .B(_6749_), .C(_6627__bF_buf3), .Y(_6757_) );
	OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf0), .B(_6342__bF_buf2), .C(_6752_), .Y(_6758_) );
	NAND3X1 NAND3X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_6757_), .C(_6758_), .Y(_6759_) );
	AOI22X1 AOI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(_6742_), .B(_6748_), .C(_6759_), .D(_6756_), .Y(_6760_) );
	XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(divider_aOp_abs_7_), .Y(_6761_) );
	INVX1 INVX1_1047 ( .gnd(gnd), .vdd(vdd), .A(_6761_), .Y(_6762_) );
	NAND3X1 NAND3X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf1), .B(_6762_), .C(_6627__bF_buf2), .Y(_6763_) );
	OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf5), .B(_6342__bF_buf1), .C(_6333_), .Y(_6764_) );
	NAND3X1 NAND3X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf0), .B(_6763_), .C(_6764_), .Y(_6765_) );
	AOI21X1 AOI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6763_), .C(_1768__bF_buf7), .Y(_6767_) );
	NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_6_), .B(_1746__bF_buf3), .Y(_6768_) );
	OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(_6767_), .C(_6765_), .Y(_6769_) );
	NAND2X1 NAND2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_6267_), .B(_6289_), .Y(_6770_) );
	INVX1 INVX1_1048 ( .gnd(gnd), .vdd(vdd), .A(_6363_), .Y(_6771_) );
	OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .B(_6771_), .C(_6362_), .Y(_6772_) );
	XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_6772_), .B(_6770_), .Y(_6773_) );
	NAND3X1 NAND3X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf0), .B(_6773_), .C(_6627__bF_buf1), .Y(_6774_) );
	OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf4), .B(_6342__bF_buf0), .C(_6266_), .Y(_6775_) );
	NAND3X1 NAND3X1_1473 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .B(_6774_), .C(_6775_), .Y(_6776_) );
	INVX1 INVX1_1049 ( .gnd(gnd), .vdd(vdd), .A(_6773_), .Y(_6778_) );
	NOR3X1 NOR3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf3), .B(_6778_), .C(_6342__bF_buf4), .Y(_6779_) );
	OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_5332__bF_buf0), .B(_5886__bF_buf1), .C(_6286_), .Y(_6780_) );
	AOI22X1 AOI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_6265_), .B(_6780_), .C(_1615__bF_buf4), .D(_6627__bF_buf0), .Y(_6781_) );
	OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_6781_), .B(_6779_), .C(_2470__bF_buf1), .Y(_6782_) );
	OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_6285_), .B(_6279_), .Y(_6783_) );
	AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_6783_), .B(_6362_), .Y(_6784_) );
	INVX1 INVX1_1050 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .Y(_6785_) );
	NAND3X1 NAND3X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf3), .B(_6785_), .C(_6627__bF_buf3), .Y(_6786_) );
	OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf2), .B(_6342__bF_buf3), .C(_6771_), .Y(_6787_) );
	NAND3X1 NAND3X1_1475 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .B(_6786_), .C(_6787_), .Y(_6789_) );
	OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf1), .B(_6342__bF_buf2), .C(_6363_), .Y(_6790_) );
	NAND3X1 NAND3X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf2), .B(_6784_), .C(_6627__bF_buf2), .Y(_6791_) );
	NAND3X1 NAND3X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_6791_), .C(_6790_), .Y(_6792_) );
	AOI22X1 AOI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(_6789_), .B(_6792_), .C(_6776_), .D(_6782_), .Y(_6793_) );
	NAND3X1 NAND3X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_6760_), .B(_6769_), .C(_6793_), .Y(_6794_) );
	NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_6735_), .B(_6794_), .Y(_6795_) );
	AOI22X1 AOI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(_6701_), .B(_6706_), .C(_6686_), .D(_6692_), .Y(_6796_) );
	AOI21X1 AOI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_6708_), .B(_6715_), .C(_4714__bF_buf3), .Y(_6797_) );
	NAND3X1 NAND3X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf2), .B(_6715_), .C(_6708_), .Y(_6798_) );
	NAND3X1 NAND3X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf0), .B(_6725_), .C(_6728_), .Y(_6800_) );
	AOI21X1 AOI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .B(_6800_), .C(_6797_), .Y(_6801_) );
	NAND3X1 NAND3X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf4), .B(_6671_), .C(_6685_), .Y(_6802_) );
	AOI21X1 AOI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_6685_), .B(_6671_), .C(_8971__bF_buf3), .Y(_6803_) );
	NAND3X1 NAND3X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf5), .B(_6698_), .C(_6699_), .Y(_6804_) );
	OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_6804_), .B(_6803_), .C(_6802_), .Y(_6805_) );
	AOI21X1 AOI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_6796_), .B(_6801_), .C(_6805_), .Y(_6806_) );
	NAND3X1 NAND3X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_6774_), .C(_6775_), .Y(_6807_) );
	AOI21X1 AOI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_6775_), .B(_6774_), .C(_2470__bF_buf7), .Y(_6808_) );
	NAND3X1 NAND3X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_6786_), .C(_6787_), .Y(_6809_) );
	OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_6809_), .B(_6808_), .C(_6807_), .Y(_6811_) );
	NAND3X1 NAND3X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf7), .B(_6741_), .C(_6736_), .Y(_6812_) );
	AOI21X1 AOI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_6736_), .B(_6741_), .C(_4100__bF_buf6), .Y(_6813_) );
	NAND3X1 NAND3X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf7), .B(_6751_), .C(_6754_), .Y(_6814_) );
	OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_6814_), .B(_6813_), .C(_6812_), .Y(_6815_) );
	AOI21X1 AOI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_6760_), .C(_6815_), .Y(_6816_) );
	OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_6735_), .B(_6816_), .C(_6806_), .Y(_6817_) );
	NAND2X1 NAND2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_6605_), .B(_6611_), .Y(_6818_) );
	NAND2X1 NAND2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_6617_), .B(_6621_), .Y(_6819_) );
	NAND3X1 NAND3X1_1487 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .B(_6624_), .C(_6640_), .Y(_6820_) );
	INVX1 INVX1_1051 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .Y(_6822_) );
	OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf0), .B(_6342__bF_buf1), .C(_6822_), .Y(_6823_) );
	NAND3X1 NAND3X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_6635_), .B(_6630_), .C(_6637_), .Y(_6824_) );
	OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_6139_), .B(_6632_), .C(_6629_), .Y(_6825_) );
	NAND2X1 NAND2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_6824_), .B(_6825_), .Y(_6826_) );
	NAND3X1 NAND3X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf1), .B(_6627__bF_buf1), .C(_6826_), .Y(_6827_) );
	NAND3X1 NAND3X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf2), .B(_6823_), .C(_6827_), .Y(_6828_) );
	NAND3X1 NAND3X1_1491 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .B(_6644_), .C(_6648_), .Y(_6829_) );
	INVX1 INVX1_1052 ( .gnd(gnd), .vdd(vdd), .A(_6643_), .Y(_6830_) );
	NAND3X1 NAND3X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_1615__bF_buf0), .B(_6830_), .C(_6627__bF_buf0), .Y(_6831_) );
	OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_4008__bF_buf5), .B(_6342__bF_buf0), .C(_6646_), .Y(_6833_) );
	NAND3X1 NAND3X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf0), .B(_6831_), .C(_6833_), .Y(_6834_) );
	AOI22X1 AOI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_6829_), .B(_6834_), .C(_6820_), .D(_6828_), .Y(_6835_) );
	NAND3X1 NAND3X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_6819_), .B(_6835_), .C(_6818_), .Y(_6836_) );
	NOR3X1 NOR3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .B(_6836_), .C(_6556_), .Y(_6837_) );
	OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_6795_), .B(_6817_), .C(_6837_), .Y(_6838_) );
	AOI21X1 AOI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_6838_), .B(_6670_), .C(_6523_), .Y(_6839_) );
	OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_6496_), .B(_6839_), .C(_6345_), .Y(_6840_) );
	AOI21X1 AOI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf6), .B(_6344_), .C(_2240__bF_buf0), .Y(_6841_) );
	INVX1 INVX1_1053 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .Y(_6842_) );
	NAND2X1 NAND2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf0), .B(_6842_), .Y(_6844_) );
	INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf3), .Y(_6845_) );
	NAND2X1 NAND2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_6841_), .Y(_6846_) );
	INVX1 INVX1_1054 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .Y(_6847_) );
	NOR3X1 NOR3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_6499_), .B(_6503_), .C(_6521_), .Y(_6848_) );
	NAND3X1 NAND3X1_1495 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf0), .B(_6525_), .C(_6537_), .Y(_6849_) );
	NAND3X1 NAND3X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf2), .B(_6540_), .C(_6543_), .Y(_6850_) );
	AOI22X1 AOI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(_6549_), .B(_6554_), .C(_6849_), .D(_6850_), .Y(_6851_) );
	NAND3X1 NAND3X1_1497 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .B(_6566_), .C(_6565_), .Y(_6852_) );
	OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_6572_), .B(_6573_), .C(_1944__bF_buf0), .Y(_6853_) );
	AOI22X1 AOI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_6580_), .B(_6584_), .C(_6852_), .D(_6853_), .Y(_6855_) );
	NAND2X1 NAND2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_6855_), .B(_6851_), .Y(_6856_) );
	AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_6662_), .B(_6574_), .Y(_6857_) );
	AOI21X1 AOI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_6537_), .B(_6525_), .C(_2887__bF_buf1), .Y(_6858_) );
	OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_6665_), .B(_6858_), .C(_6538_), .Y(_6859_) );
	AOI21X1 AOI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_6851_), .B(_6857_), .C(_6859_), .Y(_6860_) );
	OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_6657_), .B(_6856_), .C(_6860_), .Y(_6861_) );
	AOI21X1 AOI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_6848_), .B(_6861_), .C(_6496_), .Y(_6862_) );
	OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_6794_), .B(_6735_), .Y(_6863_) );
	AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_6796_), .B(_6734_), .Y(_6864_) );
	AOI21X1 AOI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_6747_), .B(_6745_), .C(_4100__bF_buf5), .Y(_6866_) );
	AOI21X1 AOI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_6736_), .B(_6741_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .Y(_6867_) );
	AOI21X1 AOI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_6758_), .B(_6757_), .C(_1735__bF_buf6), .Y(_6868_) );
	AOI21X1 AOI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_6754_), .B(_6751_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .Y(_6869_) );
	OAI22X1 OAI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_6866_), .B(_6867_), .C(_6868_), .D(_6869_), .Y(_6870_) );
	NOR3X1 NOR3X1_69 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_6781_), .C(_6779_), .Y(_6871_) );
	OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_6781_), .B(_6779_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .Y(_6872_) );
	AOI21X1 AOI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_6790_), .B(_6791_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .Y(_6873_) );
	AOI21X1 AOI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_6872_), .B(_6873_), .C(_6871_), .Y(_6874_) );
	INVX1 INVX1_1055 ( .gnd(gnd), .vdd(vdd), .A(_6812_), .Y(_6875_) );
	OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_6746_), .B(divider_divuResult_7_bF_buf5), .C(_6741_), .Y(_6877_) );
	NAND2X1 NAND2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .B(_6877_), .Y(_6878_) );
	INVX1 INVX1_1056 ( .gnd(gnd), .vdd(vdd), .A(_6814_), .Y(_6879_) );
	AOI21X1 AOI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .B(_6878_), .C(_6875_), .Y(_6880_) );
	OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_6870_), .B(_6874_), .C(_6880_), .Y(_6881_) );
	NAND2X1 NAND2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_6881_), .B(_6864_), .Y(_6882_) );
	NAND3X1 NAND3X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_6806_), .B(_6882_), .C(_6863_), .Y(_6883_) );
	NAND3X1 NAND3X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_6837_), .B(_6883_), .C(_6848_), .Y(_6884_) );
	AOI21X1 AOI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_6862_), .B(_6884_), .C(_6847_), .Y(divider_divuResult_6_) );
	NAND2X1 NAND2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_6390_), .B(_6385_), .Y(_6885_) );
	INVX1 INVX1_1057 ( .gnd(gnd), .vdd(vdd), .A(_6885_), .Y(_6887_) );
	OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_6416_), .B(divider_divuResult_7_bF_buf4), .C(_6422_), .Y(_6888_) );
	INVX1 INVX1_1058 ( .gnd(gnd), .vdd(vdd), .A(_6888_), .Y(_6889_) );
	OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf1), .B(_6889_), .C(_6486_), .Y(_6890_) );
	NAND2X1 NAND2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_6500_), .B(_6890_), .Y(_6891_) );
	NAND3X1 NAND3X1_1500 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf1), .B(_6443_), .C(_6446_), .Y(_6892_) );
	NAND3X1 NAND3X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_6481_), .B(_6892_), .C(_6506_), .Y(_6893_) );
	INVX1 INVX1_1059 ( .gnd(gnd), .vdd(vdd), .A(_6479_), .Y(_6894_) );
	INVX1 INVX1_1060 ( .gnd(gnd), .vdd(vdd), .A(_6481_), .Y(_6895_) );
	INVX1 INVX1_1061 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .Y(_6896_) );
	AOI21X1 AOI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_6892_), .B(_6896_), .C(_6895_), .Y(_6898_) );
	OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_6893_), .B(_6894_), .C(_6898_), .Y(_6899_) );
	AOI21X1 AOI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_6838_), .B(_6670_), .C(_6521_), .Y(_6900_) );
	OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_6899_), .B(_6900_), .C(_6426_), .Y(_6901_) );
	AOI21X1 AOI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_6891_), .C(_6887_), .Y(_6902_) );
	OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_6687_), .B(_6691_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .Y(_6903_) );
	NAND3X1 NAND3X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_6802_), .B(_6903_), .C(_6707_), .Y(_6904_) );
	INVX1 INVX1_1062 ( .gnd(gnd), .vdd(vdd), .A(_6797_), .Y(_6905_) );
	OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_6717_), .B(divider_divuResult_7_bF_buf3), .C(_6715_), .Y(_6906_) );
	OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .B(_6906_), .C(_6800_), .Y(_6907_) );
	NAND2X1 NAND2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_6905_), .B(_6907_), .Y(_6909_) );
	NOR3X1 NOR3X1_70 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .B(_6687_), .C(_6691_), .Y(_6910_) );
	INVX1 INVX1_1063 ( .gnd(gnd), .vdd(vdd), .A(_6804_), .Y(_6911_) );
	AOI21X1 AOI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_6911_), .B(_6903_), .C(_6910_), .Y(_6912_) );
	OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_6909_), .B(_6904_), .C(_6912_), .Y(_6913_) );
	AOI21X1 AOI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_6864_), .B(_6881_), .C(_6913_), .Y(_6914_) );
	INVX1 INVX1_1064 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .Y(_6915_) );
	NAND3X1 NAND3X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_6855_), .B(_6851_), .C(_6915_), .Y(_6916_) );
	AOI21X1 AOI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_6863_), .C(_6916_), .Y(_6917_) );
	OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6917_), .C(_6522_), .Y(_6918_) );
	AOI21X1 AOI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_6918_), .B(_6485_), .C(_6503_), .Y(_6920_) );
	NOR3X1 NOR3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_6885_), .B(_6488_), .C(_6920_), .Y(_6921_) );
	OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_6902_), .B(_6921_), .C(divider_divuResult_6_bF_buf6), .Y(_6922_) );
	NAND2X1 NAND2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_6389_), .B(_6388_), .Y(_6923_) );
	OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf5), .B(_6923_), .Y(_6924_) );
	NAND3X1 NAND3X1_1504 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_6924_), .C(_6922_), .Y(_6925_) );
	OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_6488_), .B(_6920_), .C(_6885_), .Y(_6926_) );
	NAND3X1 NAND3X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_6887_), .B(_6891_), .C(_6901_), .Y(_6927_) );
	NAND3X1 NAND3X1_1506 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf4), .B(_6927_), .C(_6926_), .Y(_6928_) );
	NAND2X1 NAND2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_6923_), .B(_6840__bF_buf5), .Y(_6929_) );
	NAND3X1 NAND3X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_6929_), .C(_6928_), .Y(_6931_) );
	AOI22X1 AOI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(_6844_), .B(_6846_), .C(_6931_), .D(_6925_), .Y(_6932_) );
	OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_6402_), .B(_6411_), .C(_6840__bF_buf4), .Y(_6933_) );
	NAND2X1 NAND2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_6401_), .B(_6412_), .Y(_6934_) );
	OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_6899_), .B(_6900_), .C(_6501_), .Y(_6935_) );
	NAND3X1 NAND3X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .B(_6418_), .C(_6935_), .Y(_6936_) );
	INVX1 INVX1_1065 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .Y(_6937_) );
	INVX1 INVX1_1066 ( .gnd(gnd), .vdd(vdd), .A(_6418_), .Y(_6938_) );
	AOI21X1 AOI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_6918_), .B(_6485_), .C(_6424_), .Y(_6939_) );
	OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6939_), .C(_6937_), .Y(_6940_) );
	NAND3X1 NAND3X1_1509 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf3), .B(_6936_), .C(_6940_), .Y(_6942_) );
	NAND3X1 NAND3X1_1510 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf1), .B(_6933_), .C(_6942_), .Y(_6943_) );
	INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(_6933_), .Y(_6944_) );
	OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6939_), .C(_6934_), .Y(_6945_) );
	NAND3X1 NAND3X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_6937_), .B(_6418_), .C(_6935_), .Y(_6946_) );
	AOI21X1 AOI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_6945_), .B(_6946_), .C(_6840__bF_buf3), .Y(_6947_) );
	OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_6944_), .B(_6947_), .C(_2042__bF_buf0), .Y(_6948_) );
	NAND3X1 NAND3X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_6424_), .B(_6485_), .C(_6918_), .Y(_6949_) );
	INVX1 INVX1_1067 ( .gnd(gnd), .vdd(vdd), .A(_6949_), .Y(_6950_) );
	OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_6939_), .B(_6950_), .C(divider_divuResult_6_bF_buf2), .Y(_6951_) );
	NAND2X1 NAND2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_6889_), .B(_6840__bF_buf2), .Y(_6953_) );
	NAND3X1 NAND3X1_1513 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf1), .B(_6953_), .C(_6951_), .Y(_6954_) );
	AOI21X1 AOI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_6949_), .B(_6935_), .C(_6840__bF_buf1), .Y(_6955_) );
	NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_6888_), .B(divider_divuResult_6_bF_buf1), .Y(_6956_) );
	OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_6956_), .B(_6955_), .C(_5516__bF_buf0), .Y(_6957_) );
	AOI22X1 AOI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_6954_), .B(_6957_), .C(_6943_), .D(_6948_), .Y(_6958_) );
	NAND2X1 NAND2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_6958_), .Y(_6959_) );
	OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_6442_), .B(divider_divuResult_7_bF_buf2), .C(_6440_), .Y(_6960_) );
	NAND2X1 NAND2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_6960_), .B(_6840__bF_buf0), .Y(_6961_) );
	INVX1 INVX1_1068 ( .gnd(gnd), .vdd(vdd), .A(_6520_), .Y(_6962_) );
	AOI21X1 AOI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_6838_), .B(_6670_), .C(_6962_), .Y(_6964_) );
	OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_6479_), .B(_6964_), .C(_6506_), .Y(_6965_) );
	NAND3X1 NAND3X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_6505_), .B(_6483_), .C(_6965_), .Y(_6966_) );
	INVX1 INVX1_1069 ( .gnd(gnd), .vdd(vdd), .A(_6505_), .Y(_6967_) );
	OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6917_), .C(_6520_), .Y(_6968_) );
	AOI22X1 AOI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(_6454_), .B(_6459_), .C(_6894_), .D(_6968_), .Y(_6969_) );
	OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6969_), .C(_6967_), .Y(_6970_) );
	NAND3X1 NAND3X1_1515 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf0), .B(_6966_), .C(_6970_), .Y(_6971_) );
	NAND3X1 NAND3X1_1516 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf0), .B(_6961_), .C(_6971_), .Y(_6972_) );
	OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_6969_), .C(_6505_), .Y(_6973_) );
	NAND3X1 NAND3X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_6967_), .B(_6483_), .C(_6965_), .Y(_6975_) );
	NAND3X1 NAND3X1_1518 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf6), .B(_6975_), .C(_6973_), .Y(_6976_) );
	INVX1 INVX1_1070 ( .gnd(gnd), .vdd(vdd), .A(_6960_), .Y(_6977_) );
	NAND2X1 NAND2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_6977_), .B(_6840__bF_buf6), .Y(_6978_) );
	NAND3X1 NAND3X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf1), .B(_6978_), .C(_6976_), .Y(_6979_) );
	AOI21X1 AOI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_6883_), .B(_6837_), .C(_6861_), .Y(_6980_) );
	OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(_6980_), .C(_6894_), .Y(_6981_) );
	NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_6506_), .B(_6981_), .Y(_6982_) );
	OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_6969_), .B(_6982_), .C(divider_divuResult_6_bF_buf5), .Y(_6983_) );
	OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_6455_), .B(_6457_), .C(_6840__bF_buf5), .Y(_6984_) );
	NAND3X1 NAND3X1_1520 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf0), .B(_6984_), .C(_6983_), .Y(_6986_) );
	NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf4), .B(_6969_), .Y(_6987_) );
	OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_6506_), .B(_6981_), .C(_6987_), .Y(_6988_) );
	OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_6456_), .B(divider_divuResult_7_bF_buf1), .C(_6452_), .Y(_6989_) );
	INVX1 INVX1_1071 ( .gnd(gnd), .vdd(vdd), .A(_6989_), .Y(_6990_) );
	NAND2X1 NAND2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_6990_), .B(_6840__bF_buf3), .Y(_6991_) );
	NAND3X1 NAND3X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf1), .B(_6991_), .C(_6988_), .Y(_6992_) );
	AOI22X1 AOI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_6986_), .B(_6992_), .C(_6972_), .D(_6979_), .Y(_6993_) );
	OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_6511_), .B(divider_divuResult_7_bF_buf0), .C(_6471_), .Y(_6994_) );
	NAND2X1 NAND2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_6994_), .B(_6840__bF_buf2), .Y(_6995_) );
	INVX1 INVX1_1072 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .Y(_6997_) );
	NAND2X1 NAND2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_6507_), .B(_6514_), .Y(_6998_) );
	AOI21X1 AOI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_6838_), .B(_6670_), .C(_6519_), .Y(_6999_) );
	OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_6997_), .B(_6999_), .C(_6998_), .Y(_7000_) );
	INVX1 INVX1_1073 ( .gnd(gnd), .vdd(vdd), .A(_6998_), .Y(_7001_) );
	INVX1 INVX1_1074 ( .gnd(gnd), .vdd(vdd), .A(_6519_), .Y(_7002_) );
	OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6917_), .C(_7002_), .Y(_7003_) );
	NAND3X1 NAND3X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .B(_7001_), .C(_7003_), .Y(_7004_) );
	NAND2X1 NAND2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_7000_), .B(_7004_), .Y(_7005_) );
	NAND2X1 NAND2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf4), .B(_7005_), .Y(_7006_) );
	NAND3X1 NAND3X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf3), .B(_6995_), .C(_7006_), .Y(_7008_) );
	NAND2X1 NAND2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_6519_), .B(_6980_), .Y(_7009_) );
	NAND2X1 NAND2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_7003_), .B(_7009_), .Y(_7010_) );
	NAND2X1 NAND2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf3), .B(_7010_), .Y(_7011_) );
	OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_6016_), .B(divider_divuResult_7_bF_buf6), .C(_6475_), .Y(_7012_) );
	NAND2X1 NAND2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_7012_), .B(_6840__bF_buf1), .Y(_7013_) );
	NAND2X1 NAND2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_7013_), .B(_7011_), .Y(_7014_) );
	INVX1 INVX1_1075 ( .gnd(gnd), .vdd(vdd), .A(_7014_), .Y(_7015_) );
	NAND2X1 NAND2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf0), .B(_7015_), .Y(_7016_) );
	AOI21X1 AOI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_7006_), .B(_6995_), .C(_4011__bF_buf2), .Y(_7017_) );
	OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_7017_), .B(_7016_), .C(_7008_), .Y(_7019_) );
	NAND3X1 NAND3X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf0), .B(_6961_), .C(_6971_), .Y(_7020_) );
	AOI21X1 AOI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_6971_), .B(_6961_), .C(_4881__bF_buf3), .Y(_7021_) );
	NAND3X1 NAND3X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf0), .B(_6984_), .C(_6983_), .Y(_7022_) );
	OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .B(_7021_), .C(_7020_), .Y(_7023_) );
	AOI21X1 AOI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_7019_), .B(_6993_), .C(_7023_), .Y(_7024_) );
	NAND3X1 NAND3X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf3), .B(_6933_), .C(_6942_), .Y(_7025_) );
	AOI21X1 AOI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_6942_), .B(_6933_), .C(_2042__bF_buf2), .Y(_7026_) );
	NAND3X1 NAND3X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf3), .B(_6953_), .C(_6951_), .Y(_7027_) );
	AOI21X1 AOI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_7027_), .C(_7026_), .Y(_7028_) );
	NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf2), .B(_6841_), .Y(_7030_) );
	INVX1 INVX1_1076 ( .gnd(gnd), .vdd(vdd), .A(_7030_), .Y(_7031_) );
	NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_6842_), .Y(_7032_) );
	NAND3X1 NAND3X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_6924_), .C(_6922_), .Y(_7033_) );
	OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_7032_), .B(_7033_), .C(_7031_), .Y(_7034_) );
	AOI21X1 AOI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_7028_), .C(_7034_), .Y(_7035_) );
	OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_6959_), .B(_7024_), .C(_7035_), .Y(_7036_) );
	NAND2X1 NAND2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_6844_), .Y(_7037_) );
	NAND3X1 NAND3X1_1529 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_6929_), .C(_6928_), .Y(_7038_) );
	NAND3X1 NAND3X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_7037_), .B(_7038_), .C(_7033_), .Y(_7039_) );
	OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_6944_), .B(_6947_), .C(divider_absoluteValue_B_flipSign_result_24_bF_buf0), .Y(_7041_) );
	NAND2X1 NAND2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_6957_), .B(_6954_), .Y(_7042_) );
	NAND3X1 NAND3X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_7042_), .C(_7041_), .Y(_7043_) );
	NAND2X1 NAND2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_6972_), .B(_6979_), .Y(_7044_) );
	NAND2X1 NAND2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_6986_), .B(_6992_), .Y(_7045_) );
	NAND3X1 NAND3X1_1532 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf2), .B(_6995_), .C(_7006_), .Y(_7046_) );
	INVX1 INVX1_1077 ( .gnd(gnd), .vdd(vdd), .A(_6994_), .Y(_7047_) );
	NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_7047_), .B(divider_divuResult_6_bF_buf2), .Y(_7048_) );
	AOI21X1 AOI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_7004_), .B(_7000_), .C(_6840__bF_buf0), .Y(_7049_) );
	OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_7048_), .B(_7049_), .C(_4011__bF_buf1), .Y(_7050_) );
	NAND3X1 NAND3X1_1533 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf2), .B(_7013_), .C(_7011_), .Y(_7052_) );
	NAND2X1 NAND2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf4), .B(_7014_), .Y(_7053_) );
	AOI22X1 AOI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(_7046_), .B(_7050_), .C(_7053_), .D(_7052_), .Y(_7054_) );
	NAND3X1 NAND3X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_7045_), .B(_7054_), .C(_7044_), .Y(_7055_) );
	NOR3X1 NOR3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_7039_), .B(_7043_), .C(_7055_), .Y(_7056_) );
	OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_6539_), .B(divider_divuResult_7_bF_buf5), .C(_6537_), .Y(_7057_) );
	NAND2X1 NAND2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_7057_), .B(_6840__bF_buf6), .Y(_7058_) );
	NAND2X1 NAND2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_6850_), .Y(_7059_) );
	OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_6795_), .B(_6817_), .C(_6915_), .Y(_7060_) );
	AOI21X1 AOI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_7060_), .B(_6657_), .C(_6586_), .Y(_7061_) );
	OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_6857_), .B(_7061_), .C(_6555_), .Y(_7063_) );
	NAND3X1 NAND3X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_7059_), .B(_6665_), .C(_7063_), .Y(_7064_) );
	INVX1 INVX1_1078 ( .gnd(gnd), .vdd(vdd), .A(_7059_), .Y(_7065_) );
	AOI21X1 AOI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_6863_), .C(_6836_), .Y(_7066_) );
	OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_7066_), .C(_6855_), .Y(_7067_) );
	AOI22X1 AOI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(_6549_), .B(_6554_), .C(_6663_), .D(_7067_), .Y(_7068_) );
	OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(_7068_), .C(_7065_), .Y(_7069_) );
	NAND3X1 NAND3X1_1536 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf1), .B(_7064_), .C(_7069_), .Y(_7070_) );
	NAND3X1 NAND3X1_1537 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf4), .B(_7058_), .C(_7070_), .Y(_7071_) );
	OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(_7068_), .C(_7059_), .Y(_7072_) );
	NAND3X1 NAND3X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_7065_), .B(_6665_), .C(_7063_), .Y(_7074_) );
	NAND3X1 NAND3X1_1539 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf0), .B(_7074_), .C(_7072_), .Y(_7075_) );
	INVX1 INVX1_1079 ( .gnd(gnd), .vdd(vdd), .A(_7057_), .Y(_7076_) );
	NAND2X1 NAND2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_7076_), .B(_6840__bF_buf5), .Y(_7077_) );
	NAND3X1 NAND3X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf3), .B(_7077_), .C(_7075_), .Y(_7078_) );
	NOR3X1 NOR3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_6555_), .B(_6857_), .C(_7061_), .Y(_7079_) );
	OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_7079_), .B(_7068_), .C(divider_divuResult_6_bF_buf6), .Y(_7080_) );
	OAI21X1 OAI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_6552_), .B(divider_divuResult_7_bF_buf4), .C(_6547_), .Y(_7081_) );
	NAND2X1 NAND2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .B(_6840__bF_buf4), .Y(_7082_) );
	NAND3X1 NAND3X1_1541 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .B(_7082_), .C(_7080_), .Y(_7083_) );
	INVX1 INVX1_1080 ( .gnd(gnd), .vdd(vdd), .A(_6555_), .Y(_7085_) );
	NAND3X1 NAND3X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_7085_), .B(_6663_), .C(_7067_), .Y(_7086_) );
	AOI21X1 AOI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_7086_), .B(_7063_), .C(_6840__bF_buf3), .Y(_7087_) );
	INVX1 INVX1_1081 ( .gnd(gnd), .vdd(vdd), .A(_7081_), .Y(_7088_) );
	NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_7088_), .B(divider_divuResult_6_bF_buf5), .Y(_7089_) );
	OAI21X1 OAI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_7089_), .B(_7087_), .C(_2887__bF_buf0), .Y(_7090_) );
	AOI22X1 AOI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(_7083_), .B(_7090_), .C(_7071_), .D(_7078_), .Y(_7091_) );
	NAND2X1 NAND2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_6852_), .B(_6853_), .Y(_7092_) );
	OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_6661_), .B(divider_absoluteValue_B_flipSign_result_14_bF_buf1), .Y(_7093_) );
	INVX1 INVX1_1082 ( .gnd(gnd), .vdd(vdd), .A(_7093_), .Y(_7094_) );
	INVX1 INVX1_1083 ( .gnd(gnd), .vdd(vdd), .A(_6585_), .Y(_7096_) );
	AOI21X1 AOI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_7060_), .B(_6657_), .C(_7096_), .Y(_7097_) );
	OAI21X1 OAI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_7094_), .B(_7097_), .C(_7092_), .Y(_7098_) );
	INVX1 INVX1_1084 ( .gnd(gnd), .vdd(vdd), .A(_7092_), .Y(_7099_) );
	OAI21X1 OAI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_7066_), .C(_6585_), .Y(_7100_) );
	NAND3X1 NAND3X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_7099_), .B(_7093_), .C(_7100_), .Y(_7101_) );
	NAND3X1 NAND3X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_7098_), .B(_7101_), .C(divider_divuResult_6_bF_buf4), .Y(_7102_) );
	NAND2X1 NAND2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_6660_), .B(_6840__bF_buf2), .Y(_7103_) );
	AOI21X1 AOI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_7102_), .B(_7103_), .C(_2922__bF_buf0), .Y(_7104_) );
	OAI21X1 OAI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_6572_), .B(_6573_), .C(_6840__bF_buf1), .Y(_7105_) );
	NAND2X1 NAND2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_7098_), .B(_7101_), .Y(_7107_) );
	NAND2X1 NAND2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf3), .B(_7107_), .Y(_7108_) );
	AOI21X1 AOI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_7108_), .B(_7105_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .Y(_7109_) );
	OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf2), .B(_6661_), .Y(_7110_) );
	NAND3X1 NAND3X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_7096_), .B(_6657_), .C(_7060_), .Y(_7111_) );
	NAND2X1 NAND2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_7111_), .B(_7100_), .Y(_7112_) );
	OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf0), .B(_7112_), .Y(_7113_) );
	AOI21X1 AOI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_7110_), .B(_7113_), .C(_1944__bF_buf4), .Y(_7114_) );
	NAND2X1 NAND2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_7112_), .B(divider_divuResult_6_bF_buf1), .Y(_7115_) );
	NAND2X1 NAND2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_6661_), .B(_6840__bF_buf6), .Y(_7116_) );
	AOI21X1 AOI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_7115_), .B(_7116_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .Y(_7118_) );
	OAI22X1 OAI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_7114_), .B(_7118_), .C(_7104_), .D(_7109_), .Y(_7119_) );
	INVX1 INVX1_1085 ( .gnd(gnd), .vdd(vdd), .A(_7119_), .Y(_7120_) );
	NAND2X1 NAND2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_7091_), .B(_7120_), .Y(_7121_) );
	OAI21X1 OAI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_6606_), .B(divider_divuResult_7_bF_buf3), .C(_6604_), .Y(_7122_) );
	NAND2X1 NAND2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_7122_), .B(_6840__bF_buf5), .Y(_7123_) );
	INVX1 INVX1_1086 ( .gnd(gnd), .vdd(vdd), .A(_6651_), .Y(_7124_) );
	OAI21X1 OAI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_6795_), .B(_6817_), .C(_6835_), .Y(_7125_) );
	AOI22X1 AOI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_6617_), .B(_6621_), .C(_7124_), .D(_7125_), .Y(_7126_) );
	INVX1 INVX1_1087 ( .gnd(gnd), .vdd(vdd), .A(_7126_), .Y(_7127_) );
	NAND3X1 NAND3X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_6818_), .B(_6654_), .C(_7127_), .Y(_7129_) );
	INVX1 INVX1_1088 ( .gnd(gnd), .vdd(vdd), .A(_6818_), .Y(_7130_) );
	INVX1 INVX1_1089 ( .gnd(gnd), .vdd(vdd), .A(_6654_), .Y(_7131_) );
	OAI21X1 OAI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_7131_), .B(_7126_), .C(_7130_), .Y(_7132_) );
	NAND3X1 NAND3X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_7132_), .B(divider_divuResult_6_bF_buf0), .C(_7129_), .Y(_7133_) );
	NAND3X1 NAND3X1_1548 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf0), .B(_7123_), .C(_7133_), .Y(_7134_) );
	INVX1 INVX1_1090 ( .gnd(gnd), .vdd(vdd), .A(_7122_), .Y(_7135_) );
	NAND2X1 NAND2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_7135_), .B(_6840__bF_buf4), .Y(_7136_) );
	OAI21X1 OAI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_7131_), .B(_7126_), .C(_6818_), .Y(_7137_) );
	NAND3X1 NAND3X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_7130_), .B(_6654_), .C(_7127_), .Y(_7138_) );
	NAND3X1 NAND3X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_7137_), .B(divider_divuResult_6_bF_buf6), .C(_7138_), .Y(_7140_) );
	NAND3X1 NAND3X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf0), .B(_7136_), .C(_7140_), .Y(_7141_) );
	NAND2X1 NAND2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(_7125_), .Y(_7142_) );
	OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_7142_), .B(_6819_), .Y(_7143_) );
	NAND2X1 NAND2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_7127_), .B(_7143_), .Y(_7144_) );
	NAND2X1 NAND2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf5), .B(_7144_), .Y(_7145_) );
	NAND3X1 NAND3X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_6619_), .B(_6620_), .C(_6840__bF_buf3), .Y(_7146_) );
	NAND3X1 NAND3X1_1553 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .B(_7146_), .C(_7145_), .Y(_7147_) );
	NAND3X1 NAND3X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_6615_), .B(_6616_), .C(_6840__bF_buf2), .Y(_7148_) );
	NAND3X1 NAND3X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_7127_), .B(_7143_), .C(divider_divuResult_6_bF_buf4), .Y(_7149_) );
	NAND3X1 NAND3X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf3), .B(_7148_), .C(_7149_), .Y(_7151_) );
	AOI22X1 AOI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_7151_), .C(_7134_), .D(_7141_), .Y(_7152_) );
	NAND2X1 NAND2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_6820_), .B(_6828_), .Y(_7153_) );
	OAI21X1 OAI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_6646_), .B(divider_divuResult_7_bF_buf2), .C(_6644_), .Y(_7154_) );
	NAND2X1 NAND2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_6829_), .B(_6834_), .Y(_7155_) );
	OAI21X1 OAI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_6795_), .B(_6817_), .C(_7155_), .Y(_7156_) );
	OAI21X1 OAI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .B(_7154_), .C(_7156_), .Y(_7157_) );
	NAND2X1 NAND2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_7153_), .B(_7157_), .Y(_7158_) );
	INVX1 INVX1_1091 ( .gnd(gnd), .vdd(vdd), .A(_7153_), .Y(_7159_) );
	NAND3X1 NAND3X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_7159_), .C(_7156_), .Y(_7160_) );
	NAND2X1 NAND2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .B(_7158_), .Y(_7162_) );
	NAND2X1 NAND2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_7162_), .B(divider_divuResult_6_bF_buf3), .Y(_7163_) );
	OAI21X1 OAI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_6408_), .B(_6826_), .C(_6624_), .Y(_7164_) );
	NAND2X1 NAND2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_7164_), .B(_6840__bF_buf1), .Y(_7165_) );
	NAND3X1 NAND3X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf4), .B(_7165_), .C(_7163_), .Y(_7166_) );
	XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_6883_), .B(_7155_), .Y(_7167_) );
	OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf0), .B(_7167_), .Y(_7168_) );
	NAND2X1 NAND2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_7154_), .B(_6840__bF_buf6), .Y(_7169_) );
	NAND3X1 NAND3X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf1), .B(_7169_), .C(_7168_), .Y(_7170_) );
	AOI21X1 AOI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_7163_), .B(_7165_), .C(_1484__bF_buf3), .Y(_7171_) );
	OAI21X1 OAI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_7171_), .B(_7170_), .C(_7166_), .Y(_7173_) );
	NAND3X1 NAND3X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf4), .B(_7123_), .C(_7133_), .Y(_7174_) );
	AOI21X1 AOI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .B(_7123_), .C(_1505__bF_buf3), .Y(_7175_) );
	NAND3X1 NAND3X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf2), .B(_7146_), .C(_7145_), .Y(_7176_) );
	OAI21X1 OAI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_7176_), .B(_7175_), .C(_7174_), .Y(_7177_) );
	AOI21X1 AOI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_7152_), .B(_7173_), .C(_7177_), .Y(_7178_) );
	AOI21X1 AOI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_7102_), .B(_7103_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf4), .Y(_7179_) );
	INVX1 INVX1_1092 ( .gnd(gnd), .vdd(vdd), .A(_7179_), .Y(_7180_) );
	AOI21X1 AOI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_7108_), .B(_7105_), .C(_2922__bF_buf3), .Y(_7181_) );
	AOI21X1 AOI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_7110_), .B(_7113_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .Y(_7182_) );
	INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(_7182_), .Y(_7184_) );
	AOI21X1 AOI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_7184_), .B(_7180_), .C(_7181_), .Y(_7185_) );
	NAND3X1 NAND3X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf2), .B(_7058_), .C(_7070_), .Y(_7186_) );
	AOI21X1 AOI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_7070_), .B(_7058_), .C(_3263__bF_buf1), .Y(_7187_) );
	OAI21X1 OAI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_7088_), .B(divider_divuResult_6_bF_buf2), .C(_7080_), .Y(_7188_) );
	OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_7188_), .B(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .Y(_7189_) );
	OAI21X1 OAI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_7187_), .B(_7189_), .C(_7186_), .Y(_7190_) );
	AOI21X1 AOI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_7185_), .B(_7091_), .C(_7190_), .Y(_7191_) );
	OAI21X1 OAI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_7178_), .B(_7121_), .C(_7191_), .Y(_7192_) );
	AOI21X1 AOI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_7056_), .B(_7192_), .C(_7036_), .Y(_7193_) );
	INVX1 INVX1_1093 ( .gnd(gnd), .vdd(vdd), .A(_6734_), .Y(_7194_) );
	AOI21X1 AOI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_6816_), .B(_6794_), .C(_7194_), .Y(_7195_) );
	OAI21X1 OAI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_6801_), .B(_7195_), .C(_6707_), .Y(_7196_) );
	NAND3X1 NAND3X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_6693_), .B(_6804_), .C(_7196_), .Y(_7197_) );
	INVX1 INVX1_1094 ( .gnd(gnd), .vdd(vdd), .A(_6707_), .Y(_7198_) );
	NAND2X1 NAND2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_6794_), .B(_6816_), .Y(_7199_) );
	AOI21X1 AOI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_7199_), .B(_6734_), .C(_6801_), .Y(_7200_) );
	OAI21X1 OAI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_7198_), .B(_7200_), .C(_6804_), .Y(_7201_) );
	OAI21X1 OAI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_6910_), .B(_6803_), .C(_7201_), .Y(_7202_) );
	NAND2X1 NAND2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_7197_), .B(_7202_), .Y(_7203_) );
	OAI21X1 OAI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_6687_), .B(_6691_), .C(_6840__bF_buf5), .Y(_7205_) );
	OAI21X1 OAI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf4), .B(_7203_), .C(_7205_), .Y(_7206_) );
	NAND2X1 NAND2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .B(_7206_), .Y(_7207_) );
	NAND2X1 NAND2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_6693_), .B(_7201_), .Y(_7208_) );
	INVX1 INVX1_1095 ( .gnd(gnd), .vdd(vdd), .A(_6693_), .Y(_7209_) );
	NAND3X1 NAND3X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_7209_), .B(_6804_), .C(_7196_), .Y(_7210_) );
	NAND2X1 NAND2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_7210_), .B(_7208_), .Y(_7211_) );
	NAND2X1 NAND2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_7211_), .B(divider_divuResult_6_bF_buf1), .Y(_7212_) );
	NAND3X1 NAND3X1_1565 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .B(_7205_), .C(_7212_), .Y(_7213_) );
	NAND2X1 NAND2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_7203_), .B(divider_divuResult_6_bF_buf0), .Y(_7214_) );
	OAI21X1 OAI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_6214_), .B(divider_divuResult_7_bF_buf1), .C(_6685_), .Y(_7216_) );
	INVX1 INVX1_1096 ( .gnd(gnd), .vdd(vdd), .A(_7216_), .Y(_7217_) );
	NAND2X1 NAND2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_7217_), .B(_6840__bF_buf3), .Y(_7218_) );
	NAND3X1 NAND3X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf5), .B(_7218_), .C(_7214_), .Y(_7219_) );
	AOI21X1 AOI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_6388_), .B(_6389_), .C(divider_absoluteValue_B_flipSign_result_24_bF_buf3), .Y(_7220_) );
	AOI21X1 AOI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_7220_), .B(_6497_), .C(_6489_), .Y(_7221_) );
	OAI21X1 OAI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_6499_), .B(_6891_), .C(_7221_), .Y(_7222_) );
	AOI21X1 AOI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_6899_), .B(_6504_), .C(_7222_), .Y(_7223_) );
	NAND2X1 NAND2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_6848_), .B(_6861_), .Y(_7224_) );
	NAND3X1 NAND3X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_7223_), .B(_7224_), .C(_6884_), .Y(_7225_) );
	NAND2X1 NAND2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_7198_), .B(_7200_), .Y(_7227_) );
	NAND2X1 NAND2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_7196_), .B(_7227_), .Y(_7228_) );
	NAND3X1 NAND3X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7228_), .C(_7225_), .Y(_7229_) );
	OAI21X1 OAI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(divider_divuResult_7_bF_buf0), .C(_6698_), .Y(_7230_) );
	NAND2X1 NAND2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7230_), .B(_6840__bF_buf2), .Y(_7231_) );
	NAND3X1 NAND3X1_1569 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .B(_7229_), .C(_7231_), .Y(_7232_) );
	INVX1 INVX1_1097 ( .gnd(gnd), .vdd(vdd), .A(_7228_), .Y(_7233_) );
	NAND3X1 NAND3X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7225_), .C(_7233_), .Y(_7234_) );
	INVX1 INVX1_1098 ( .gnd(gnd), .vdd(vdd), .A(_7230_), .Y(_7235_) );
	NAND2X1 NAND2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_7235_), .B(_6840__bF_buf1), .Y(_7236_) );
	NAND3X1 NAND3X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf2), .B(_7234_), .C(_7236_), .Y(_7238_) );
	AOI22X1 AOI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(_7232_), .B(_7238_), .C(_7213_), .D(_7219_), .Y(_7239_) );
	NAND3X1 NAND3X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf4), .B(_7205_), .C(_7212_), .Y(_7240_) );
	OAI21X1 OAI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_7235_), .B(divider_divuResult_6_bF_buf6), .C(_7229_), .Y(_7241_) );
	OAI21X1 OAI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .B(_7241_), .C(_7240_), .Y(_7242_) );
	NAND2X1 NAND2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_6906_), .B(_6840__bF_buf0), .Y(_7243_) );
	NAND2X1 NAND2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_6716_), .B(_6721_), .Y(_7244_) );
	OAI21X1 OAI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_6726_), .B(divider_divuResult_7_bF_buf6), .C(_6725_), .Y(_7245_) );
	NAND2X1 NAND2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_6729_), .B(_6732_), .Y(_7246_) );
	NAND2X1 NAND2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_7246_), .B(_7199_), .Y(_7247_) );
	OAI21X1 OAI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_7245_), .C(_7247_), .Y(_7249_) );
	XNOR2X1 XNOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_7249_), .B(_7244_), .Y(_7250_) );
	NAND3X1 NAND3X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7225_), .C(_7250_), .Y(_7251_) );
	AOI21X1 AOI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_7243_), .B(_7251_), .C(_7204__bF_buf4), .Y(_7252_) );
	NAND3X1 NAND3X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_7251_), .C(_7243_), .Y(_7253_) );
	XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_7199_), .B(_7246_), .Y(_7254_) );
	INVX1 INVX1_1099 ( .gnd(gnd), .vdd(vdd), .A(_7254_), .Y(_7255_) );
	NAND3X1 NAND3X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7255_), .C(_7225_), .Y(_7256_) );
	NAND2X1 NAND2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_7245_), .B(_6840__bF_buf6), .Y(_7257_) );
	NAND3X1 NAND3X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf1), .B(_7256_), .C(_7257_), .Y(_7258_) );
	AOI21X1 AOI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_7253_), .B(_7258_), .C(_7252_), .Y(_7260_) );
	AOI22X1 AOI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(_7207_), .B(_7242_), .C(_7260_), .D(_7239_), .Y(_7261_) );
	NAND3X1 NAND3X1_1577 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_7251_), .C(_7243_), .Y(_7262_) );
	INVX1 INVX1_1100 ( .gnd(gnd), .vdd(vdd), .A(_6906_), .Y(_7263_) );
	NAND2X1 NAND2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_7263_), .B(_6840__bF_buf5), .Y(_7264_) );
	XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_7249_), .B(_7244_), .Y(_7265_) );
	NAND3X1 NAND3X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7225_), .C(_7265_), .Y(_7266_) );
	NAND3X1 NAND3X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf2), .B(_7266_), .C(_7264_), .Y(_7267_) );
	NAND3X1 NAND3X1_1580 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .B(_7256_), .C(_7257_), .Y(_7268_) );
	NAND3X1 NAND3X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_6725_), .B(_6728_), .C(_6840__bF_buf4), .Y(_7269_) );
	NAND2X1 NAND2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_7254_), .B(divider_divuResult_6_bF_buf5), .Y(_7271_) );
	NAND3X1 NAND3X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf0), .B(_7269_), .C(_7271_), .Y(_7272_) );
	AOI22X1 AOI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(_7262_), .B(_7267_), .C(_7268_), .D(_7272_), .Y(_7273_) );
	AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_7273_), .B(_7239_), .Y(_7274_) );
	INVX1 INVX1_1101 ( .gnd(gnd), .vdd(vdd), .A(_6765_), .Y(_7275_) );
	NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_6767_), .B(_7275_), .Y(_7276_) );
	XNOR2X1 XNOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_7276_), .B(_6768_), .Y(_7277_) );
	NAND3X1 NAND3X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7277_), .C(_7225_), .Y(_7278_) );
	NAND3X1 NAND3X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_6763_), .B(_6764_), .C(_6840__bF_buf3), .Y(_7279_) );
	NAND3X1 NAND3X1_1585 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_7278_), .C(_7279_), .Y(_7280_) );
	INVX1 INVX1_1102 ( .gnd(gnd), .vdd(vdd), .A(_7280_), .Y(_7282_) );
	OAI21X1 OAI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_7_), .B(divider_divuResult_7_bF_buf5), .C(_6763_), .Y(_7283_) );
	OAI21X1 OAI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_7283_), .B(divider_divuResult_6_bF_buf4), .C(_7278_), .Y(_7284_) );
	INVX1 INVX1_1103 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_6_), .Y(_7285_) );
	XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(divider_aOp_abs_6_), .Y(_7286_) );
	INVX1 INVX1_1104 ( .gnd(gnd), .vdd(vdd), .A(_7286_), .Y(_7287_) );
	MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_7285_), .B(_7287_), .S(_6840__bF_buf2), .Y(_7288_) );
	AOI22X1 AOI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(_7284_), .B(_2547__bF_buf1), .C(_1768__bF_buf6), .D(_7288_), .Y(_7289_) );
	NAND2X1 NAND2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_7287_), .B(divider_divuResult_6_bF_buf3), .Y(_7290_) );
	NAND2X1 NAND2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_7285_), .B(_6840__bF_buf1), .Y(_7291_) );
	NAND3X1 NAND3X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_7291_), .C(_7290_), .Y(_7293_) );
	OAI21X1 OAI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf2), .B(_6840__bF_buf0), .C(divider_aOp_abs_6_), .Y(_7294_) );
	NAND2X1 NAND2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(divider_divuResult_6_bF_buf2), .Y(_7295_) );
	NAND3X1 NAND3X1_1587 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .B(_7295_), .C(_7294_), .Y(_7296_) );
	NAND2X1 NAND2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_7293_), .B(_7296_), .Y(_7297_) );
	INVX1 INVX1_1105 ( .gnd(gnd), .vdd(vdd), .A(_7277_), .Y(_7298_) );
	NAND3X1 NAND3X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7298_), .C(_7225_), .Y(_7299_) );
	NAND2X1 NAND2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_7283_), .B(_6840__bF_buf6), .Y(_7300_) );
	NAND3X1 NAND3X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf0), .B(_7299_), .C(_7300_), .Y(_7301_) );
	NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_5_), .B(_1746__bF_buf1), .Y(_7302_) );
	INVX1 INVX1_1106 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .Y(_7304_) );
	NAND3X1 NAND3X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_7304_), .B(_7301_), .C(_7280_), .Y(_7305_) );
	OAI22X1 OAI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_7282_), .B(_7289_), .C(_7305_), .D(_7297_), .Y(_7306_) );
	NAND2X1 NAND2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .B(_6840__bF_buf5), .Y(_7307_) );
	NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_6866_), .B(_6867_), .Y(_7308_) );
	NAND2X1 NAND2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_6759_), .Y(_7309_) );
	INVX1 INVX1_1107 ( .gnd(gnd), .vdd(vdd), .A(_6769_), .Y(_7310_) );
	INVX1 INVX1_1108 ( .gnd(gnd), .vdd(vdd), .A(_6793_), .Y(_7311_) );
	OAI21X1 OAI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_7310_), .B(_7311_), .C(_6874_), .Y(_7312_) );
	AOI21X1 AOI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_7309_), .C(_6879_), .Y(_7313_) );
	XNOR2X1 XNOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_7313_), .B(_7308_), .Y(_7315_) );
	NAND3X1 NAND3X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7315_), .C(_7225_), .Y(_7316_) );
	NAND3X1 NAND3X1_1592 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_7316_), .C(_7307_), .Y(_7317_) );
	INVX1 INVX1_1109 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .Y(_7318_) );
	OAI21X1 OAI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_7318_), .B(divider_divuResult_6_bF_buf1), .C(_7316_), .Y(_7319_) );
	NAND2X1 NAND2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf6), .B(_7319_), .Y(_7320_) );
	XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_7309_), .Y(_7321_) );
	INVX1 INVX1_1110 ( .gnd(gnd), .vdd(vdd), .A(_7321_), .Y(_7322_) );
	NAND3X1 NAND3X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7322_), .C(_7225_), .Y(_7323_) );
	OAI21X1 OAI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_6752_), .B(divider_divuResult_7_bF_buf4), .C(_6751_), .Y(_7324_) );
	NAND2X1 NAND2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_7324_), .B(_6840__bF_buf4), .Y(_7326_) );
	NAND3X1 NAND3X1_1594 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_7323_), .C(_7326_), .Y(_7327_) );
	NAND3X1 NAND3X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7321_), .C(_7225_), .Y(_7328_) );
	INVX1 INVX1_1111 ( .gnd(gnd), .vdd(vdd), .A(_7324_), .Y(_7329_) );
	NAND2X1 NAND2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(_6840__bF_buf3), .Y(_7330_) );
	NAND3X1 NAND3X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf4), .B(_7328_), .C(_7330_), .Y(_7331_) );
	AOI22X1 AOI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(_7327_), .B(_7331_), .C(_7317_), .D(_7320_), .Y(_7332_) );
	NAND2X1 NAND2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_6776_), .B(_6782_), .Y(_7333_) );
	INVX1 INVX1_1112 ( .gnd(gnd), .vdd(vdd), .A(_6789_), .Y(_7334_) );
	INVX1 INVX1_1113 ( .gnd(gnd), .vdd(vdd), .A(_6792_), .Y(_7335_) );
	NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_7334_), .B(_7335_), .Y(_7337_) );
	OAI21X1 OAI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_7337_), .B(_7310_), .C(_6809_), .Y(_7338_) );
	XNOR2X1 XNOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_7338_), .B(_7333_), .Y(_7339_) );
	NAND3X1 NAND3X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7339_), .C(_7225_), .Y(_7340_) );
	OAI21X1 OAI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_6779_), .B(_6781_), .C(_6840__bF_buf2), .Y(_7341_) );
	NAND3X1 NAND3X1_1598 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .B(_7340_), .C(_7341_), .Y(_7342_) );
	OAI21X1 OAI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_6288_), .B(divider_divuResult_7_bF_buf3), .C(_6774_), .Y(_7343_) );
	INVX1 INVX1_1114 ( .gnd(gnd), .vdd(vdd), .A(_7343_), .Y(_7344_) );
	OAI21X1 OAI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_7344_), .B(divider_divuResult_6_bF_buf0), .C(_7340_), .Y(_7345_) );
	NAND2X1 NAND2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf5), .B(_7345_), .Y(_7346_) );
	XNOR2X1 XNOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_7337_), .B(_6769_), .Y(_7348_) );
	INVX1 INVX1_1115 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .Y(_7349_) );
	NAND3X1 NAND3X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7349_), .C(_7225_), .Y(_7350_) );
	OAI21X1 OAI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_6363_), .B(divider_divuResult_7_bF_buf2), .C(_6786_), .Y(_7351_) );
	NAND2X1 NAND2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .B(_6840__bF_buf1), .Y(_7352_) );
	NAND3X1 NAND3X1_1600 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .B(_7350_), .C(_7352_), .Y(_7353_) );
	NAND3X1 NAND3X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_6345_), .B(_7348_), .C(_7225_), .Y(_7354_) );
	INVX1 INVX1_1116 ( .gnd(gnd), .vdd(vdd), .A(_7351_), .Y(_7355_) );
	NAND2X1 NAND2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_7355_), .B(_6840__bF_buf0), .Y(_7356_) );
	NAND3X1 NAND3X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_7354_), .C(_7356_), .Y(_7357_) );
	AOI22X1 AOI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(_7353_), .B(_7357_), .C(_7342_), .D(_7346_), .Y(_7359_) );
	AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7359_), .Y(_7360_) );
	NAND3X1 NAND3X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_7306_), .B(_7274_), .C(_7360_), .Y(_7361_) );
	NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_7319_), .Y(_7362_) );
	AOI21X1 AOI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .B(_7316_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .Y(_7363_) );
	AOI21X1 AOI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_7330_), .B(_7328_), .C(_4100__bF_buf3), .Y(_7364_) );
	AOI21X1 AOI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_7326_), .B(_7323_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .Y(_7365_) );
	OAI22X1 OAI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_7364_), .B(_7365_), .C(_7363_), .D(_7362_), .Y(_7366_) );
	NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .B(_7345_), .Y(_7367_) );
	NAND2X1 NAND2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_7345_), .Y(_7368_) );
	AOI21X1 AOI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_7356_), .B(_7354_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .Y(_7370_) );
	AOI21X1 AOI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_7368_), .B(_7370_), .C(_7367_), .Y(_7371_) );
	NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_7319_), .Y(_7372_) );
	NAND2X1 NAND2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .B(_7319_), .Y(_7373_) );
	NAND3X1 NAND3X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_7323_), .C(_7326_), .Y(_7374_) );
	INVX1 INVX1_1117 ( .gnd(gnd), .vdd(vdd), .A(_7374_), .Y(_7375_) );
	AOI21X1 AOI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_7373_), .C(_7372_), .Y(_7376_) );
	OAI21X1 OAI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_7371_), .B(_7366_), .C(_7376_), .Y(_7377_) );
	NAND2X1 NAND2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_7274_), .B(_7377_), .Y(_7378_) );
	NAND3X1 NAND3X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_7261_), .B(_7361_), .C(_7378_), .Y(_7379_) );
	NAND3X1 NAND3X1_1606 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf3), .B(_7077_), .C(_7075_), .Y(_7381_) );
	NAND2X1 NAND2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_7083_), .B(_7090_), .Y(_7382_) );
	NAND3X1 NAND3X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_7186_), .C(_7381_), .Y(_7383_) );
	NAND3X1 NAND3X1_1608 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .B(_7165_), .C(_7163_), .Y(_7384_) );
	AOI21X1 AOI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_7158_), .B(_7160_), .C(_6840__bF_buf6), .Y(_7385_) );
	AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf5), .B(_7164_), .Y(_7386_) );
	OAI21X1 OAI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_7385_), .B(_7386_), .C(_1484__bF_buf2), .Y(_7387_) );
	NAND3X1 NAND3X1_1609 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .B(_7169_), .C(_7168_), .Y(_7388_) );
	NAND2X1 NAND2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .B(divider_divuResult_6_bF_buf6), .Y(_7389_) );
	NAND3X1 NAND3X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_6648_), .C(_6840__bF_buf4), .Y(_7390_) );
	NAND3X1 NAND3X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf0), .B(_7390_), .C(_7389_), .Y(_7392_) );
	AOI22X1 AOI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7392_), .C(_7384_), .D(_7387_), .Y(_7393_) );
	NAND2X1 NAND2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7152_), .Y(_7394_) );
	NOR3X1 NOR3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_7119_), .B(_7383_), .C(_7394_), .Y(_7395_) );
	NAND3X1 NAND3X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_7395_), .B(_7056_), .C(_7379_), .Y(_7396_) );
	AOI21X1 AOI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_7193_), .B(_7396_), .C(_6315__bF_buf4), .Y(divider_divuResult_5_) );
	NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_7119_), .B(_7383_), .Y(_7397_) );
	AOI21X1 AOI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_7140_), .B(_7136_), .C(_1505__bF_buf2), .Y(_7398_) );
	AOI21X1 AOI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .B(_7123_), .C(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .Y(_7399_) );
	AOI21X1 AOI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_7149_), .B(_7148_), .C(_1494__bF_buf1), .Y(_7400_) );
	AOI21X1 AOI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_7145_), .B(_7146_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .Y(_7402_) );
	OAI22X1 OAI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_7402_), .C(_7398_), .D(_7399_), .Y(_7403_) );
	INVX1 INVX1_1118 ( .gnd(gnd), .vdd(vdd), .A(_7166_), .Y(_7404_) );
	AOI21X1 AOI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_7389_), .B(_7390_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .Y(_7405_) );
	OAI21X1 OAI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_7385_), .B(_7386_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .Y(_7406_) );
	AOI21X1 AOI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_7406_), .C(_7404_), .Y(_7407_) );
	INVX1 INVX1_1119 ( .gnd(gnd), .vdd(vdd), .A(_7174_), .Y(_7408_) );
	NAND3X1 NAND3X1_1613 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .B(_7136_), .C(_7140_), .Y(_7409_) );
	AOI21X1 AOI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_7149_), .B(_7148_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .Y(_7410_) );
	AOI21X1 AOI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_7410_), .B(_7409_), .C(_7408_), .Y(_7411_) );
	OAI21X1 OAI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_7407_), .B(_7403_), .C(_7411_), .Y(_7413_) );
	OAI21X1 OAI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_6660_), .B(divider_divuResult_6_bF_buf5), .C(_7108_), .Y(_7414_) );
	NAND2X1 NAND2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf3), .B(_7414_), .Y(_7415_) );
	OAI21X1 OAI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_7179_), .B(_7182_), .C(_7415_), .Y(_7416_) );
	AOI21X1 AOI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_7075_), .B(_7077_), .C(divider_absoluteValue_B_flipSign_result_18_bF_buf2), .Y(_7417_) );
	NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .B(_7188_), .Y(_7418_) );
	AOI21X1 AOI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_7381_), .B(_7418_), .C(_7417_), .Y(_7419_) );
	OAI21X1 OAI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_7416_), .B(_7383_), .C(_7419_), .Y(_7420_) );
	AOI21X1 AOI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_7397_), .B(_7413_), .C(_7420_), .Y(_7421_) );
	NAND2X1 NAND2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_7239_), .B(_7273_), .Y(_7422_) );
	NAND2X1 NAND2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_7422_), .B(_7261_), .Y(_7424_) );
	OAI21X1 OAI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf3), .B(_7277_), .C(_7300_), .Y(_7425_) );
	OAI21X1 OAI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .B(_7425_), .C(_7293_), .Y(_7426_) );
	OAI21X1 OAI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_7284_), .C(_7426_), .Y(_7427_) );
	NAND3X1 NAND3X1_1614 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .B(_7291_), .C(_7290_), .Y(_7428_) );
	NAND3X1 NAND3X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_7295_), .C(_7294_), .Y(_7429_) );
	NAND2X1 NAND2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .B(_7429_), .Y(_7430_) );
	INVX1 INVX1_1120 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_5_), .Y(_7431_) );
	NAND3X1 NAND3X1_1616 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_7299_), .C(_7300_), .Y(_7432_) );
	NAND3X1 NAND3X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf6), .B(_7278_), .C(_7279_), .Y(_7433_) );
	AOI22X1 AOI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(_7431_), .C(_7432_), .D(_7433_), .Y(_7435_) );
	NAND2X1 NAND2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_7430_), .B(_7435_), .Y(_7436_) );
	NAND2X1 NAND2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7359_), .Y(_7437_) );
	AOI21X1 AOI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_7427_), .B(_7436_), .C(_7437_), .Y(_7438_) );
	NAND3X1 NAND3X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf4), .B(_7340_), .C(_7341_), .Y(_7439_) );
	AOI21X1 AOI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_7341_), .B(_7340_), .C(_1735__bF_buf3), .Y(_7440_) );
	NAND3X1 NAND3X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf5), .B(_7350_), .C(_7352_), .Y(_7441_) );
	OAI21X1 OAI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_7441_), .B(_7440_), .C(_7439_), .Y(_7442_) );
	NAND2X1 NAND2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_7442_), .B(_7332_), .Y(_7443_) );
	NAND3X1 NAND3X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_7376_), .B(_7443_), .C(_7261_), .Y(_7444_) );
	OAI21X1 OAI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_7438_), .B(_7444_), .C(_7424_), .Y(_7446_) );
	AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_7152_), .B(_7393_), .Y(_7447_) );
	NAND3X1 NAND3X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_7091_), .B(_7120_), .C(_7447_), .Y(_7448_) );
	OAI21X1 OAI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_7448_), .B(_7446_), .C(_7421_), .Y(_7449_) );
	AOI21X1 AOI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_7449_), .B(_7056_), .C(_7036_), .Y(_7450_) );
	OAI21X1 OAI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_6842_), .Y(_7451_) );
	AOI21X1 AOI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_7451_), .B(_2229__bF_buf2), .C(divider_absoluteValue_B_flipSign_result_27_), .Y(_7452_) );
	INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .Y(_7453_) );
	OAI21X1 OAI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(divider_divuResult_5_bF_buf6), .C(_2229__bF_buf1), .Y(_7454_) );
	NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_7454_), .Y(_7455_) );
	NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_7452_), .B(_7455_), .Y(_7457_) );
	NAND2X1 NAND2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .B(_6925_), .Y(_7458_) );
	INVX1 INVX1_1121 ( .gnd(gnd), .vdd(vdd), .A(_7458_), .Y(_7459_) );
	NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_6944_), .B(_6947_), .Y(_7460_) );
	OAI21X1 OAI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_6888_), .B(divider_divuResult_6_bF_buf4), .C(_6951_), .Y(_7461_) );
	OAI21X1 OAI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf0), .B(_7461_), .C(_7025_), .Y(_7462_) );
	OAI21X1 OAI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf1), .B(_7460_), .C(_7462_), .Y(_7463_) );
	NAND2X1 NAND2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_7045_), .B(_7044_), .Y(_7464_) );
	OAI21X1 OAI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_7047_), .B(divider_divuResult_6_bF_buf3), .C(_7006_), .Y(_7465_) );
	INVX1 INVX1_1122 ( .gnd(gnd), .vdd(vdd), .A(_7465_), .Y(_7466_) );
	OAI21X1 OAI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf1), .B(_7014_), .C(_7008_), .Y(_7468_) );
	OAI21X1 OAI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf0), .B(_7466_), .C(_7468_), .Y(_7469_) );
	INVX1 INVX1_1123 ( .gnd(gnd), .vdd(vdd), .A(_7020_), .Y(_7470_) );
	OAI21X1 OAI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_6977_), .B(divider_divuResult_6_bF_buf2), .C(_6971_), .Y(_7471_) );
	NAND2X1 NAND2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf3), .B(_7471_), .Y(_7472_) );
	INVX1 INVX1_1124 ( .gnd(gnd), .vdd(vdd), .A(_7022_), .Y(_7473_) );
	AOI21X1 AOI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_7472_), .B(_7473_), .C(_7470_), .Y(_7474_) );
	OAI21X1 OAI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_7469_), .B(_7464_), .C(_7474_), .Y(_7475_) );
	AOI22X1 AOI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(_7426_), .B(_7280_), .C(_7430_), .D(_7435_), .Y(_7476_) );
	NOR3X1 NOR3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_7422_), .B(_7437_), .C(_7476_), .Y(_7477_) );
	MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .B(_7315_), .S(_6840__bF_buf2), .Y(_7479_) );
	NAND2X1 NAND2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_7479_), .Y(_7480_) );
	AOI21X1 AOI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_7307_), .B(_7316_), .C(_4999__bF_buf3), .Y(_7481_) );
	OAI21X1 OAI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .B(_7374_), .C(_7480_), .Y(_7482_) );
	AOI21X1 AOI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7442_), .C(_7482_), .Y(_7483_) );
	OAI21X1 OAI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_7422_), .B(_7483_), .C(_7261_), .Y(_7484_) );
	OAI21X1 OAI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_7484_), .B(_7477_), .C(_7395_), .Y(_7485_) );
	AOI21X1 AOI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .B(_7421_), .C(_7055_), .Y(_7486_) );
	OAI21X1 OAI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_7475_), .B(_7486_), .C(_6958_), .Y(_7487_) );
	AOI21X1 AOI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_7487_), .B(_7463_), .C(_7459_), .Y(_7488_) );
	NAND3X1 NAND3X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_7459_), .B(_7463_), .C(_7487_), .Y(_7490_) );
	INVX1 INVX1_1125 ( .gnd(gnd), .vdd(vdd), .A(_7490_), .Y(_7491_) );
	OAI21X1 OAI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_7488_), .B(_7491_), .C(divider_divuResult_5_bF_buf5), .Y(_7492_) );
	NAND2X1 NAND2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_6929_), .B(_6928_), .Y(_7493_) );
	OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf4), .B(_7493_), .Y(_7494_) );
	NAND3X1 NAND3X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_7494_), .C(_7492_), .Y(_7495_) );
	INVX1 INVX1_1126 ( .gnd(gnd), .vdd(vdd), .A(_7055_), .Y(_7496_) );
	AOI21X1 AOI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_7449_), .B(_7496_), .C(_7475_), .Y(_7497_) );
	OAI21X1 OAI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_7043_), .B(_7497_), .C(_7463_), .Y(_7498_) );
	NAND2X1 NAND2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_7458_), .B(_7498_), .Y(_7499_) );
	NAND3X1 NAND3X1_1624 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf3), .B(_7490_), .C(_7499_), .Y(_7501_) );
	OAI21X1 OAI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(_7493_), .Y(_7502_) );
	NAND3X1 NAND3X1_1625 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf1), .B(_7502_), .C(_7501_), .Y(_7503_) );
	NAND3X1 NAND3X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_7457_), .B(_7503_), .C(_7495_), .Y(_7504_) );
	NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_7039_), .B(_7043_), .Y(_7505_) );
	NAND2X1 NAND2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_7496_), .B(_7505_), .Y(_7506_) );
	AOI21X1 AOI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .B(_7421_), .C(_7506_), .Y(_7507_) );
	OAI21X1 OAI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_7036_), .B(_7507_), .C(_6314_), .Y(_7508_) );
	OAI21X1 OAI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_6944_), .B(_6947_), .C(_7508_), .Y(_7509_) );
	NAND2X1 NAND2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_6948_), .Y(_7510_) );
	OAI21X1 OAI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_7475_), .B(_7486_), .C(_7042_), .Y(_7512_) );
	NAND3X1 NAND3X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_7510_), .B(_7027_), .C(_7512_), .Y(_7513_) );
	INVX1 INVX1_1127 ( .gnd(gnd), .vdd(vdd), .A(_7510_), .Y(_7514_) );
	INVX1 INVX1_1128 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .Y(_7515_) );
	INVX1 INVX1_1129 ( .gnd(gnd), .vdd(vdd), .A(_7206_), .Y(_7516_) );
	OAI21X1 OAI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf3), .B(_7516_), .C(_7242_), .Y(_7517_) );
	NAND2X1 NAND2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(_7239_), .Y(_7518_) );
	NAND2X1 NAND2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_7517_), .B(_7518_), .Y(_7519_) );
	AOI21X1 AOI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_7377_), .B(_7274_), .C(_7519_), .Y(_7520_) );
	AOI21X1 AOI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_7520_), .B(_7361_), .C(_7448_), .Y(_7521_) );
	OAI21X1 OAI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .B(_7521_), .C(_7496_), .Y(_7523_) );
	AOI22X1 AOI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(_6954_), .B(_6957_), .C(_7024_), .D(_7523_), .Y(_7524_) );
	OAI21X1 OAI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_7515_), .B(_7524_), .C(_7514_), .Y(_7525_) );
	NAND3X1 NAND3X1_1628 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf2), .B(_7513_), .C(_7525_), .Y(_7526_) );
	NAND3X1 NAND3X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_7509_), .C(_7526_), .Y(_7527_) );
	INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(_7509_), .Y(_7528_) );
	OAI21X1 OAI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_7515_), .B(_7524_), .C(_7510_), .Y(_7529_) );
	NAND3X1 NAND3X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_7514_), .B(_7027_), .C(_7512_), .Y(_7530_) );
	AOI21X1 AOI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_7529_), .B(_7530_), .C(_7508_), .Y(_7531_) );
	OAI21X1 OAI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_7528_), .B(_7531_), .C(divider_absoluteValue_B_flipSign_result_25_), .Y(_7532_) );
	NOR3X1 NOR3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_7042_), .B(_7475_), .C(_7486_), .Y(_7534_) );
	OAI21X1 OAI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_7524_), .B(_7534_), .C(divider_divuResult_5_bF_buf1), .Y(_7535_) );
	OAI21X1 OAI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7461_), .Y(_7536_) );
	NAND3X1 NAND3X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf0), .B(_7536_), .C(_7535_), .Y(_7537_) );
	INVX1 INVX1_1130 ( .gnd(gnd), .vdd(vdd), .A(_7042_), .Y(_7538_) );
	NAND2X1 NAND2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_7538_), .B(_7497_), .Y(_7539_) );
	NAND3X1 NAND3X1_1632 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf0), .B(_7512_), .C(_7539_), .Y(_7540_) );
	NAND3X1 NAND3X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_6951_), .B(_6953_), .C(_7508_), .Y(_7541_) );
	NAND3X1 NAND3X1_1634 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf2), .B(_7541_), .C(_7540_), .Y(_7542_) );
	AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_7537_), .B(_7542_), .Y(_7543_) );
	NAND3X1 NAND3X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_7527_), .B(_7543_), .C(_7532_), .Y(_7545_) );
	NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_7545_), .B(_7504_), .Y(_7546_) );
	OAI21X1 OAI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7471_), .Y(_7547_) );
	INVX1 INVX1_1131 ( .gnd(gnd), .vdd(vdd), .A(_7054_), .Y(_7548_) );
	AOI21X1 AOI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .B(_7421_), .C(_7548_), .Y(_7549_) );
	OAI21X1 OAI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_7019_), .B(_7549_), .C(_7045_), .Y(_7550_) );
	NAND3X1 NAND3X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_7044_), .B(_7022_), .C(_7550_), .Y(_7551_) );
	INVX1 INVX1_1132 ( .gnd(gnd), .vdd(vdd), .A(_7044_), .Y(_7552_) );
	INVX1 INVX1_1133 ( .gnd(gnd), .vdd(vdd), .A(_7045_), .Y(_7553_) );
	OAI21X1 OAI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .B(_7521_), .C(_7054_), .Y(_7554_) );
	AOI21X1 AOI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_7554_), .B(_7469_), .C(_7553_), .Y(_7556_) );
	OAI21X1 OAI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7556_), .C(_7552_), .Y(_7557_) );
	NAND3X1 NAND3X1_1637 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf6), .B(_7551_), .C(_7557_), .Y(_7558_) );
	NAND3X1 NAND3X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf2), .B(_7547_), .C(_7558_), .Y(_7559_) );
	INVX1 INVX1_1134 ( .gnd(gnd), .vdd(vdd), .A(_7471_), .Y(_7560_) );
	OAI21X1 OAI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7560_), .Y(_7561_) );
	OAI21X1 OAI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_7473_), .B(_7556_), .C(_7044_), .Y(_7562_) );
	NAND3X1 NAND3X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_7552_), .B(_7022_), .C(_7550_), .Y(_7563_) );
	NAND3X1 NAND3X1_1640 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf5), .B(_7563_), .C(_7562_), .Y(_7564_) );
	NAND3X1 NAND3X1_1641 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf3), .B(_7561_), .C(_7564_), .Y(_7565_) );
	NOR3X1 NOR3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_7045_), .B(_7019_), .C(_7549_), .Y(_7567_) );
	OAI21X1 OAI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_7567_), .B(_7556_), .C(divider_divuResult_5_bF_buf4), .Y(_7568_) );
	OAI21X1 OAI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_6990_), .B(divider_divuResult_6_bF_buf1), .C(_6983_), .Y(_7569_) );
	OAI21X1 OAI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf4), .B(_7450__bF_buf0), .C(_7569_), .Y(_7570_) );
	NAND3X1 NAND3X1_1642 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf2), .B(_7570_), .C(_7568_), .Y(_7571_) );
	NAND3X1 NAND3X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_7553_), .B(_7469_), .C(_7554_), .Y(_7572_) );
	AOI21X1 AOI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_7572_), .B(_7550_), .C(_7508_), .Y(_7573_) );
	INVX1 INVX1_1135 ( .gnd(gnd), .vdd(vdd), .A(_7569_), .Y(_7574_) );
	NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_7574_), .B(divider_divuResult_5_bF_buf3), .Y(_7575_) );
	OAI21X1 OAI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_7575_), .B(_7573_), .C(_4881__bF_buf2), .Y(_7576_) );
	NAND2X1 NAND2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_7576_), .B(_7571_), .Y(_7578_) );
	NAND3X1 NAND3X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_7578_), .B(_7559_), .C(_7565_), .Y(_7579_) );
	INVX1 INVX1_1136 ( .gnd(gnd), .vdd(vdd), .A(_7016_), .Y(_7580_) );
	NAND2X1 NAND2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_7050_), .B(_7046_), .Y(_7581_) );
	INVX1 INVX1_1137 ( .gnd(gnd), .vdd(vdd), .A(_7581_), .Y(_7582_) );
	NAND2X1 NAND2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_7052_), .B(_7053_), .Y(_7583_) );
	INVX1 INVX1_1138 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .Y(_7584_) );
	AOI21X1 AOI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_7379_), .B(_7395_), .C(_7192_), .Y(_7585_) );
	NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .B(_7585_), .Y(_7586_) );
	OAI21X1 OAI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_7580_), .B(_7586_), .C(_7582_), .Y(_7587_) );
	OAI21X1 OAI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_7192_), .B(_7521_), .C(_7583_), .Y(_7589_) );
	NAND3X1 NAND3X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_7016_), .B(_7581_), .C(_7589_), .Y(_7590_) );
	NAND3X1 NAND3X1_1646 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf2), .B(_7590_), .C(_7587_), .Y(_7591_) );
	OAI21X1 OAI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_7466_), .B(divider_divuResult_5_bF_buf1), .C(_7591_), .Y(_7592_) );
	INVX1 INVX1_1139 ( .gnd(gnd), .vdd(vdd), .A(_7592_), .Y(_7593_) );
	NAND2X1 NAND2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_7584_), .B(_7585_), .Y(_7594_) );
	NAND2X1 NAND2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_7594_), .Y(_7595_) );
	OAI21X1 OAI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_7015_), .Y(_7596_) );
	OAI21X1 OAI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7595_), .C(_7596_), .Y(_7597_) );
	NAND2X1 NAND2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf3), .B(_7597_), .Y(_7598_) );
	OAI21X1 OAI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf3), .B(_7592_), .C(_7598_), .Y(_7600_) );
	OAI21X1 OAI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf3), .B(_7593_), .C(_7600_), .Y(_7601_) );
	AOI21X1 AOI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_7564_), .B(_7561_), .C(divider_absoluteValue_B_flipSign_result_23_bF_buf2), .Y(_7602_) );
	OAI21X1 OAI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_7574_), .B(divider_divuResult_5_bF_buf0), .C(_7568_), .Y(_7603_) );
	NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf1), .B(_7603_), .Y(_7604_) );
	AOI21X1 AOI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_7565_), .B(_7604_), .C(_7602_), .Y(_7605_) );
	OAI21X1 OAI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_7579_), .B(_7601_), .C(_7605_), .Y(_7606_) );
	NOR3X1 NOR3X1_78 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_7528_), .C(_7531_), .Y(_7607_) );
	INVX1 INVX1_1140 ( .gnd(gnd), .vdd(vdd), .A(_7537_), .Y(_7608_) );
	AOI21X1 AOI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_7532_), .B(_7608_), .C(_7607_), .Y(_7609_) );
	AOI21X1 AOI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_7501_), .B(_7502_), .C(divider_absoluteValue_B_flipSign_result_26_bF_buf0), .Y(_7611_) );
	AOI21X1 AOI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_7611_), .B(_7457_), .C(_7452_), .Y(_7612_) );
	OAI21X1 OAI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_7504_), .B(_7609_), .C(_7612_), .Y(_7613_) );
	AOI21X1 AOI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_7546_), .B(_7606_), .C(_7613_), .Y(_7614_) );
	INVX1 INVX1_1141 ( .gnd(gnd), .vdd(vdd), .A(_7457_), .Y(_7615_) );
	NAND3X1 NAND3X1_1647 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf3), .B(_7494_), .C(_7492_), .Y(_7616_) );
	NAND3X1 NAND3X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_7502_), .C(_7501_), .Y(_7617_) );
	AOI21X1 AOI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_7616_), .B(_7617_), .C(_7615_), .Y(_7618_) );
	NAND3X1 NAND3X1_1649 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_7509_), .C(_7526_), .Y(_7619_) );
	OAI21X1 OAI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_7528_), .B(_7531_), .C(_2053_), .Y(_7620_) );
	NAND2X1 NAND2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_7542_), .B(_7537_), .Y(_7622_) );
	AOI21X1 AOI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_7620_), .B(_7619_), .C(_7622_), .Y(_7623_) );
	NAND2X1 NAND2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_7623_), .B(_7618_), .Y(_7624_) );
	AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_7565_), .B(_7559_), .Y(_7625_) );
	OAI21X1 OAI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(_7465_), .Y(_7626_) );
	NAND3X1 NAND3X1_1650 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf2), .B(_7626_), .C(_7591_), .Y(_7627_) );
	OAI21X1 OAI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_7580_), .B(_7586_), .C(_7581_), .Y(_7628_) );
	NAND3X1 NAND3X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_7016_), .B(_7582_), .C(_7589_), .Y(_7629_) );
	NAND3X1 NAND3X1_1652 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf6), .B(_7629_), .C(_7628_), .Y(_7630_) );
	OAI21X1 OAI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7466_), .Y(_7631_) );
	NAND3X1 NAND3X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf2), .B(_7631_), .C(_7630_), .Y(_7633_) );
	NAND2X1 NAND2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_7627_), .B(_7633_), .Y(_7634_) );
	XNOR2X1 XNOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_7597_), .B(divider_absoluteValue_B_flipSign_result_20_bF_buf1), .Y(_7635_) );
	AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .B(_7635_), .Y(_7636_) );
	NAND3X1 NAND3X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_7578_), .B(_7625_), .C(_7636_), .Y(_7637_) );
	NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_7637_), .B(_7624_), .Y(_7638_) );
	OAI21X1 OAI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_7076_), .B(divider_divuResult_6_bF_buf0), .C(_7070_), .Y(_7639_) );
	OAI21X1 OAI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7639_), .Y(_7640_) );
	NAND2X1 NAND2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_7071_), .B(_7078_), .Y(_7641_) );
	OAI21X1 OAI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_7484_), .B(_7477_), .C(_7447_), .Y(_7642_) );
	AOI21X1 AOI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_7642_), .B(_7178_), .C(_7119_), .Y(_7644_) );
	OAI21X1 OAI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_7185_), .B(_7644_), .C(_7382_), .Y(_7645_) );
	NAND3X1 NAND3X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_7641_), .B(_7189_), .C(_7645_), .Y(_7646_) );
	INVX1 INVX1_1142 ( .gnd(gnd), .vdd(vdd), .A(_7641_), .Y(_7647_) );
	INVX1 INVX1_1143 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .Y(_7648_) );
	OAI21X1 OAI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_7394_), .B(_7446_), .C(_7178_), .Y(_7649_) );
	NAND2X1 NAND2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_7120_), .B(_7649_), .Y(_7650_) );
	AOI21X1 AOI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_7650_), .B(_7416_), .C(_7648_), .Y(_7651_) );
	OAI21X1 OAI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_7418_), .B(_7651_), .C(_7647_), .Y(_7652_) );
	NAND3X1 NAND3X1_1656 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf5), .B(_7646_), .C(_7652_), .Y(_7653_) );
	NAND3X1 NAND3X1_1657 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf0), .B(_7640_), .C(_7653_), .Y(_7655_) );
	OAI21X1 OAI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_7418_), .B(_7651_), .C(_7641_), .Y(_7656_) );
	NAND3X1 NAND3X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_7647_), .B(_7189_), .C(_7645_), .Y(_7657_) );
	NAND3X1 NAND3X1_1659 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf4), .B(_7657_), .C(_7656_), .Y(_7658_) );
	INVX1 INVX1_1144 ( .gnd(gnd), .vdd(vdd), .A(_7639_), .Y(_7659_) );
	OAI21X1 OAI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7659_), .Y(_7660_) );
	NAND3X1 NAND3X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf3), .B(_7660_), .C(_7658_), .Y(_7661_) );
	NOR3X1 NOR3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_7185_), .C(_7644_), .Y(_7662_) );
	OAI21X1 OAI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(_7651_), .C(divider_divuResult_5_bF_buf3), .Y(_7663_) );
	OAI21X1 OAI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf4), .B(_7450__bF_buf0), .C(_7188_), .Y(_7664_) );
	NAND3X1 NAND3X1_1661 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf1), .B(_7664_), .C(_7663_), .Y(_7666_) );
	NAND3X1 NAND3X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_7648_), .B(_7416_), .C(_7650_), .Y(_7667_) );
	AOI21X1 AOI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_7667_), .B(_7645_), .C(_7508_), .Y(_7668_) );
	INVX1 INVX1_1145 ( .gnd(gnd), .vdd(vdd), .A(_7188_), .Y(_7669_) );
	NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_7669_), .B(divider_divuResult_5_bF_buf2), .Y(_7670_) );
	OAI21X1 OAI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_7670_), .B(_7668_), .C(_3263__bF_buf0), .Y(_7671_) );
	AOI22X1 AOI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(_7666_), .B(_7671_), .C(_7655_), .D(_7661_), .Y(_7672_) );
	INVX1 INVX1_1146 ( .gnd(gnd), .vdd(vdd), .A(_7414_), .Y(_7673_) );
	OAI21X1 OAI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_7673_), .Y(_7674_) );
	NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .B(_7114_), .Y(_7675_) );
	AOI21X1 AOI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_7379_), .B(_7447_), .C(_7413_), .Y(_7677_) );
	OAI21X1 OAI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_7675_), .B(_7677_), .C(_7184_), .Y(_7678_) );
	OAI21X1 OAI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_7104_), .B(_7109_), .C(_7678_), .Y(_7679_) );
	NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_7179_), .B(_7181_), .Y(_7680_) );
	INVX1 INVX1_1147 ( .gnd(gnd), .vdd(vdd), .A(_7680_), .Y(_7681_) );
	OAI21X1 OAI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_7114_), .B(_7118_), .C(_7649_), .Y(_7682_) );
	NAND3X1 NAND3X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_7681_), .B(_7184_), .C(_7682_), .Y(_7683_) );
	NAND3X1 NAND3X1_1664 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf1), .B(_7683_), .C(_7679_), .Y(_7684_) );
	AOI21X1 AOI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_7684_), .B(_7674_), .C(_2887__bF_buf4), .Y(_7685_) );
	INVX1 INVX1_1148 ( .gnd(gnd), .vdd(vdd), .A(_7685_), .Y(_7686_) );
	NAND3X1 NAND3X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf3), .B(_7674_), .C(_7684_), .Y(_7688_) );
	NAND2X1 NAND2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_7675_), .B(_7677_), .Y(_7689_) );
	NAND2X1 NAND2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_7682_), .B(_7689_), .Y(_7690_) );
	OAI21X1 OAI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_6661_), .B(divider_divuResult_6_bF_buf6), .C(_7113_), .Y(_7691_) );
	OAI21X1 OAI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(_7691_), .Y(_7692_) );
	OAI21X1 OAI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7690_), .C(_7692_), .Y(_7693_) );
	AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_7693_), .B(divider_absoluteValue_B_flipSign_result_16_bF_buf2), .Y(_7694_) );
	INVX1 INVX1_1149 ( .gnd(gnd), .vdd(vdd), .A(_7694_), .Y(_7695_) );
	NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf1), .B(_7693_), .Y(_7696_) );
	INVX1 INVX1_1150 ( .gnd(gnd), .vdd(vdd), .A(_7696_), .Y(_7697_) );
	AOI22X1 AOI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(_7695_), .B(_7697_), .C(_7686_), .D(_7688_), .Y(_7699_) );
	NAND2X1 NAND2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_7672_), .B(_7699_), .Y(_7700_) );
	OAI21X1 OAI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_7135_), .B(divider_divuResult_6_bF_buf5), .C(_7133_), .Y(_7701_) );
	OAI21X1 OAI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7701_), .Y(_7702_) );
	NAND2X1 NAND2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_7134_), .B(_7141_), .Y(_7703_) );
	INVX1 INVX1_1151 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .Y(_7704_) );
	OAI21X1 OAI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_7704_), .B(_7446_), .C(_7407_), .Y(_7705_) );
	OAI21X1 OAI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_7402_), .C(_7705_), .Y(_7706_) );
	NAND3X1 NAND3X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_7703_), .B(_7176_), .C(_7706_), .Y(_7707_) );
	INVX1 INVX1_1152 ( .gnd(gnd), .vdd(vdd), .A(_7703_), .Y(_7708_) );
	NAND2X1 NAND2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_7151_), .B(_7147_), .Y(_7710_) );
	INVX1 INVX1_1153 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .Y(_7711_) );
	OAI21X1 OAI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_7484_), .B(_7477_), .C(_7393_), .Y(_7712_) );
	AOI21X1 AOI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_7712_), .B(_7407_), .C(_7711_), .Y(_7713_) );
	OAI21X1 OAI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_7410_), .B(_7713_), .C(_7708_), .Y(_7714_) );
	NAND3X1 NAND3X1_1667 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf0), .B(_7714_), .C(_7707_), .Y(_7715_) );
	NAND3X1 NAND3X1_1668 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .B(_7702_), .C(_7715_), .Y(_7716_) );
	INVX1 INVX1_1154 ( .gnd(gnd), .vdd(vdd), .A(_7701_), .Y(_7717_) );
	OAI21X1 OAI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7717_), .Y(_7718_) );
	OAI21X1 OAI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_7410_), .B(_7713_), .C(_7703_), .Y(_7719_) );
	NAND3X1 NAND3X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_7708_), .B(_7176_), .C(_7706_), .Y(_7721_) );
	NAND3X1 NAND3X1_1670 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf6), .B(_7719_), .C(_7721_), .Y(_7722_) );
	NAND3X1 NAND3X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf3), .B(_7718_), .C(_7722_), .Y(_7723_) );
	AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_7716_), .B(_7723_), .Y(_7724_) );
	NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .B(_7705_), .Y(_7725_) );
	OAI21X1 OAI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_7713_), .B(_7725_), .C(divider_divuResult_5_bF_buf5), .Y(_7726_) );
	NAND3X1 NAND3X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_7148_), .B(_7149_), .C(_7508_), .Y(_7727_) );
	NAND3X1 NAND3X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf1), .B(_7726_), .C(_7727_), .Y(_7728_) );
	OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_7705_), .B(_7710_), .Y(_7729_) );
	NAND3X1 NAND3X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_7706_), .B(_7729_), .C(divider_divuResult_5_bF_buf4), .Y(_7730_) );
	OAI21X1 OAI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf1), .B(_7144_), .C(_7148_), .Y(_7732_) );
	OAI21X1 OAI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7732_), .Y(_7733_) );
	NAND3X1 NAND3X1_1675 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .B(_7733_), .C(_7730_), .Y(_7734_) );
	NAND2X1 NAND2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_7734_), .B(_7728_), .Y(_7735_) );
	NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_7735_), .B(_7724_), .Y(_7736_) );
	NAND2X1 NAND2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_7384_), .B(_7387_), .Y(_7737_) );
	NAND2X1 NAND2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_7392_), .B(_7388_), .Y(_7738_) );
	OAI21X1 OAI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_7484_), .B(_7477_), .C(_7738_), .Y(_7739_) );
	INVX1 INVX1_1155 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .Y(_7740_) );
	OAI21X1 OAI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_7740_), .C(_7737_), .Y(_7741_) );
	INVX1 INVX1_1156 ( .gnd(gnd), .vdd(vdd), .A(_7737_), .Y(_7743_) );
	NAND3X1 NAND3X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_7170_), .B(_7743_), .C(_7739_), .Y(_7744_) );
	NAND2X1 NAND2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_7744_), .B(_7741_), .Y(_7745_) );
	NAND2X1 NAND2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf3), .B(_7745_), .Y(_7746_) );
	OAI21X1 OAI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_7385_), .B(_7386_), .C(_7508_), .Y(_7747_) );
	NAND3X1 NAND3X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf0), .B(_7747_), .C(_7746_), .Y(_7748_) );
	OAI21X1 OAI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_7154_), .B(divider_divuResult_6_bF_buf4), .C(_7389_), .Y(_7749_) );
	INVX1 INVX1_1157 ( .gnd(gnd), .vdd(vdd), .A(_7749_), .Y(_7750_) );
	NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_7738_), .B(_7379_), .Y(_7751_) );
	NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_7751_), .B(_7740_), .Y(_7752_) );
	NAND2X1 NAND2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_7752_), .B(divider_divuResult_5_bF_buf2), .Y(_7754_) );
	OAI21X1 OAI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_7750_), .B(divider_divuResult_5_bF_buf1), .C(_7754_), .Y(_7755_) );
	NAND2X1 NAND2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf1), .B(_7755_), .Y(_7756_) );
	AOI21X1 AOI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .B(_7747_), .C(_1494__bF_buf4), .Y(_7757_) );
	OAI21X1 OAI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_7757_), .B(_7756_), .C(_7748_), .Y(_7758_) );
	OAI21X1 OAI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_7717_), .B(divider_divuResult_5_bF_buf0), .C(_7715_), .Y(_7759_) );
	NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .B(_7759_), .Y(_7760_) );
	INVX1 INVX1_1158 ( .gnd(gnd), .vdd(vdd), .A(_7760_), .Y(_7761_) );
	OAI21X1 OAI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .B(_7724_), .C(_7761_), .Y(_7762_) );
	AOI21X1 AOI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_7736_), .B(_7758_), .C(_7762_), .Y(_7763_) );
	AOI21X1 AOI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_7684_), .B(_7674_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .Y(_7765_) );
	INVX1 INVX1_1159 ( .gnd(gnd), .vdd(vdd), .A(_7765_), .Y(_7766_) );
	OAI21X1 OAI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf4), .B(_7450__bF_buf0), .C(_7414_), .Y(_7767_) );
	AOI21X1 AOI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_7682_), .B(_7184_), .C(_7681_), .Y(_7768_) );
	NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_7680_), .B(_7678_), .Y(_7769_) );
	OAI21X1 OAI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_7768_), .B(_7769_), .C(divider_divuResult_5_bF_buf6), .Y(_7770_) );
	AOI21X1 AOI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_7770_), .B(_7767_), .C(_2887__bF_buf2), .Y(_7771_) );
	NAND2X1 NAND2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf2), .B(_7693_), .Y(_7772_) );
	AOI21X1 AOI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_7766_), .B(_7772_), .C(_7771_), .Y(_7773_) );
	NAND3X1 NAND3X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf2), .B(_7640_), .C(_7653_), .Y(_7774_) );
	AOI21X1 AOI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_7653_), .B(_7640_), .C(_3789__bF_buf1), .Y(_7776_) );
	OAI21X1 OAI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_7669_), .B(divider_divuResult_5_bF_buf5), .C(_7663_), .Y(_7777_) );
	OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_7777_), .B(divider_absoluteValue_B_flipSign_result_18_bF_buf0), .Y(_7778_) );
	OAI21X1 OAI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_7776_), .B(_7778_), .C(_7774_), .Y(_7779_) );
	AOI21X1 AOI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_7672_), .B(_7773_), .C(_7779_), .Y(_7780_) );
	OAI21X1 OAI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_7700_), .B(_7763_), .C(_7780_), .Y(_7781_) );
	NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf0), .B(_7431_), .Y(_7782_) );
	NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7782_), .Y(_7783_) );
	AOI21X1 AOI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_6928_), .B(_6929_), .C(divider_absoluteValue_B_flipSign_result_25_), .Y(_7784_) );
	AOI21X1 AOI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_7784_), .B(_7037_), .C(_7030_), .Y(_7785_) );
	OAI21X1 OAI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_7039_), .B(_7463_), .C(_7785_), .Y(_7787_) );
	AOI21X1 AOI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_7475_), .B(_7505_), .C(_7787_), .Y(_7788_) );
	NOR3X1 NOR3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_7383_), .B(_7119_), .C(_7178_), .Y(_7789_) );
	OAI21X1 OAI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_7420_), .B(_7789_), .C(_7056_), .Y(_7790_) );
	NAND3X1 NAND3X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_7788_), .B(_7790_), .C(_7396_), .Y(_7791_) );
	NAND3X1 NAND3X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7783_), .C(_7791_), .Y(_7792_) );
	OAI21X1 OAI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_7431_), .Y(_7793_) );
	NAND3X1 NAND3X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_7792_), .C(_7793_), .Y(_7794_) );
	INVX1 INVX1_1160 ( .gnd(gnd), .vdd(vdd), .A(_7783_), .Y(_7795_) );
	NAND3X1 NAND3X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7795_), .C(_7791_), .Y(_7796_) );
	OAI21X1 OAI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(divider_aOp_abs_5_), .Y(_7797_) );
	NAND3X1 NAND3X1_1683 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .B(_7796_), .C(_7797_), .Y(_7798_) );
	AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_7794_), .B(_7798_), .Y(_7799_) );
	NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_4_), .B(_1746__bF_buf0), .Y(_7800_) );
	INVX1 INVX1_1161 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_4_), .Y(_7801_) );
	NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf5), .B(_7801_), .Y(_7802_) );
	NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_7800_), .B(_7802_), .Y(_7803_) );
	NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7297_), .Y(_7804_) );
	INVX1 INVX1_1162 ( .gnd(gnd), .vdd(vdd), .A(_7804_), .Y(_7805_) );
	NAND2X1 NAND2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7297_), .Y(_7806_) );
	NAND2X1 NAND2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_7805_), .Y(_7809_) );
	NAND3X1 NAND3X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7809_), .C(_7791_), .Y(_7810_) );
	INVX1 INVX1_1163 ( .gnd(gnd), .vdd(vdd), .A(_7288_), .Y(_7811_) );
	OAI21X1 OAI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7811_), .Y(_7812_) );
	NAND3X1 NAND3X1_1685 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_7810_), .C(_7812_), .Y(_7813_) );
	OAI21X1 OAI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7288_), .Y(_7814_) );
	INVX1 INVX1_1164 ( .gnd(gnd), .vdd(vdd), .A(_7809_), .Y(_7815_) );
	NAND3X1 NAND3X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7815_), .C(_7791_), .Y(_7816_) );
	NAND3X1 NAND3X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_7816_), .C(_7814_), .Y(_7817_) );
	OAI21X1 OAI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7425_), .Y(_7818_) );
	NAND2X1 NAND2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_7432_), .B(_7433_), .Y(_7820_) );
	OAI21X1 OAI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .B(_7297_), .C(_7293_), .Y(_7821_) );
	XNOR2X1 XNOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_7821_), .B(_7820_), .Y(_7822_) );
	NAND2X1 NAND2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_7822_), .B(divider_divuResult_5_bF_buf4), .Y(_7823_) );
	NAND3X1 NAND3X1_1688 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .B(_7818_), .C(_7823_), .Y(_7824_) );
	INVX1 INVX1_1165 ( .gnd(gnd), .vdd(vdd), .A(_7822_), .Y(_7825_) );
	NAND2X1 NAND2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_7825_), .B(divider_divuResult_5_bF_buf3), .Y(_7826_) );
	OAI21X1 OAI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf4), .B(_7450__bF_buf0), .C(_7284_), .Y(_7827_) );
	NAND3X1 NAND3X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf4), .B(_7827_), .C(_7826_), .Y(_7828_) );
	AOI22X1 AOI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .B(_7817_), .C(_7824_), .D(_7828_), .Y(_7829_) );
	NAND3X1 NAND3X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_7803_), .B(_7799_), .C(_7829_), .Y(_7831_) );
	NAND3X1 NAND3X1_1691 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .B(_7827_), .C(_7826_), .Y(_7832_) );
	AOI21X1 AOI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_7814_), .B(_7816_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .Y(_7833_) );
	AOI21X1 AOI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_7826_), .B(_7827_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .Y(_7834_) );
	AOI21X1 AOI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_7833_), .B(_7832_), .C(_7834_), .Y(_7835_) );
	AOI21X1 AOI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_7793_), .B(_7792_), .C(_1768__bF_buf2), .Y(_7836_) );
	INVX1 INVX1_1166 ( .gnd(gnd), .vdd(vdd), .A(_7802_), .Y(_7837_) );
	OAI21X1 OAI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_7837_), .B(_7836_), .C(_7794_), .Y(_7838_) );
	NAND2X1 NAND2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_7829_), .B(_7838_), .Y(_7839_) );
	NAND3X1 NAND3X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_7835_), .B(_7839_), .C(_7831_), .Y(_7840_) );
	OAI21X1 OAI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_7206_), .Y(_7842_) );
	NAND2X1 NAND2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_7219_), .B(_7213_), .Y(_7843_) );
	NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .B(_7241_), .Y(_7844_) );
	INVX1 INVX1_1167 ( .gnd(gnd), .vdd(vdd), .A(_7844_), .Y(_7845_) );
	NAND2X1 NAND2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_7232_), .B(_7238_), .Y(_7846_) );
	INVX1 INVX1_1168 ( .gnd(gnd), .vdd(vdd), .A(_7846_), .Y(_7847_) );
	OAI21X1 OAI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_7437_), .B(_7476_), .C(_7483_), .Y(_7848_) );
	AOI21X1 AOI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_7848_), .B(_7273_), .C(_7260_), .Y(_7849_) );
	OAI21X1 OAI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_7847_), .B(_7849_), .C(_7845_), .Y(_7850_) );
	AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_7850_), .B(_7843_), .Y(_7851_) );
	NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_7843_), .B(_7850_), .Y(_7853_) );
	OAI21X1 OAI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_7853_), .B(_7851_), .C(divider_divuResult_5_bF_buf2), .Y(_7854_) );
	NAND3X1 NAND3X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_7842_), .C(_7854_), .Y(_7855_) );
	NAND2X1 NAND2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_7843_), .B(_7850_), .Y(_7856_) );
	OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_7850_), .B(_7843_), .Y(_7857_) );
	NAND3X1 NAND3X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_7856_), .B(_7857_), .C(divider_divuResult_5_bF_buf1), .Y(_7858_) );
	OAI21X1 OAI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(_7516_), .Y(_7859_) );
	NAND3X1 NAND3X1_1695 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .B(_7859_), .C(_7858_), .Y(_7860_) );
	XNOR2X1 XNOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_7849_), .B(_7847_), .Y(_7861_) );
	NAND3X1 NAND3X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7861_), .C(_7791_), .Y(_7862_) );
	OAI21X1 OAI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7241_), .Y(_7864_) );
	NAND3X1 NAND3X1_1697 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .B(_7862_), .C(_7864_), .Y(_7865_) );
	XNOR2X1 XNOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_7849_), .B(_7846_), .Y(_7866_) );
	NAND3X1 NAND3X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7866_), .C(_7791_), .Y(_7867_) );
	INVX1 INVX1_1169 ( .gnd(gnd), .vdd(vdd), .A(_7241_), .Y(_7868_) );
	OAI21X1 OAI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7868_), .Y(_7869_) );
	NAND3X1 NAND3X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf2), .B(_7867_), .C(_7869_), .Y(_7870_) );
	NAND2X1 NAND2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_7865_), .B(_7870_), .Y(_7871_) );
	NAND3X1 NAND3X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_7855_), .B(_7860_), .C(_7871_), .Y(_7872_) );
	OAI21X1 OAI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_7263_), .B(divider_divuResult_6_bF_buf3), .C(_7251_), .Y(_7873_) );
	OAI21X1 OAI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7873_), .Y(_7875_) );
	NAND2X1 NAND2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_7262_), .B(_7267_), .Y(_7876_) );
	OAI21X1 OAI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_6840__bF_buf0), .B(_7254_), .C(_7257_), .Y(_7877_) );
	NAND2X1 NAND2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_7268_), .B(_7272_), .Y(_7878_) );
	OAI21X1 OAI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_7377_), .B(_7438_), .C(_7878_), .Y(_7879_) );
	OAI21X1 OAI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_7877_), .C(_7879_), .Y(_7880_) );
	NAND2X1 NAND2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_7876_), .B(_7880_), .Y(_7881_) );
	INVX1 INVX1_1170 ( .gnd(gnd), .vdd(vdd), .A(_7876_), .Y(_7882_) );
	NAND3X1 NAND3X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_7882_), .B(_7258_), .C(_7879_), .Y(_7883_) );
	NAND2X1 NAND2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_7883_), .B(_7881_), .Y(_7884_) );
	NAND3X1 NAND3X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7791_), .C(_7884_), .Y(_7886_) );
	NAND3X1 NAND3X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf1), .B(_7886_), .C(_7875_), .Y(_7887_) );
	INVX1 INVX1_1171 ( .gnd(gnd), .vdd(vdd), .A(_7873_), .Y(_7888_) );
	OAI21X1 OAI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf4), .B(_7450__bF_buf0), .C(_7888_), .Y(_7889_) );
	NAND3X1 NAND3X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_7876_), .B(_7258_), .C(_7879_), .Y(_7890_) );
	NAND2X1 NAND2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_7882_), .B(_7880_), .Y(_7891_) );
	NAND2X1 NAND2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_7890_), .B(_7891_), .Y(_7892_) );
	NAND2X1 NAND2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_7892_), .B(divider_divuResult_5_bF_buf0), .Y(_7893_) );
	NAND3X1 NAND3X1_1705 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .B(_7889_), .C(_7893_), .Y(_7894_) );
	OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_7848_), .B(_7878_), .Y(_7895_) );
	NAND2X1 NAND2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_7879_), .B(_7895_), .Y(_7897_) );
	NAND2X1 NAND2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_7897_), .B(divider_divuResult_5_bF_buf6), .Y(_7898_) );
	OAI21X1 OAI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_7877_), .Y(_7899_) );
	NAND3X1 NAND3X1_1706 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_7899_), .C(_7898_), .Y(_7900_) );
	INVX1 INVX1_1172 ( .gnd(gnd), .vdd(vdd), .A(_7877_), .Y(_7901_) );
	OAI21X1 OAI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(_7901_), .Y(_7902_) );
	INVX1 INVX1_1173 ( .gnd(gnd), .vdd(vdd), .A(_7897_), .Y(_7903_) );
	NAND2X1 NAND2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_7903_), .B(divider_divuResult_5_bF_buf5), .Y(_7904_) );
	NAND3X1 NAND3X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf1), .B(_7902_), .C(_7904_), .Y(_7905_) );
	NAND2X1 NAND2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .B(_7905_), .Y(_7906_) );
	NAND3X1 NAND3X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_7887_), .B(_7894_), .C(_7906_), .Y(_7908_) );
	NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_7872_), .B(_7908_), .Y(_7909_) );
	OAI21X1 OAI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7319_), .Y(_7910_) );
	NAND2X1 NAND2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_7317_), .B(_7320_), .Y(_7911_) );
	NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_7364_), .B(_7365_), .Y(_7912_) );
	AOI21X1 AOI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_7306_), .B(_7359_), .C(_7442_), .Y(_7913_) );
	OAI21X1 OAI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_7912_), .B(_7913_), .C(_7374_), .Y(_7914_) );
	XNOR2X1 XNOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_7914_), .B(_7911_), .Y(_7915_) );
	NAND3X1 NAND3X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7915_), .C(_7791_), .Y(_7916_) );
	NAND3X1 NAND3X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf6), .B(_7916_), .C(_7910_), .Y(_7917_) );
	OAI21X1 OAI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_7479_), .B(divider_divuResult_5_bF_buf4), .C(_7916_), .Y(_7919_) );
	NAND2X1 NAND2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .B(_7919_), .Y(_7920_) );
	XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_7913_), .B(_7912_), .Y(_7921_) );
	INVX1 INVX1_1174 ( .gnd(gnd), .vdd(vdd), .A(_7921_), .Y(_7922_) );
	NAND3X1 NAND3X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7922_), .C(_7791_), .Y(_7923_) );
	OAI21X1 OAI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .B(divider_divuResult_6_bF_buf2), .C(_7323_), .Y(_7924_) );
	OAI21X1 OAI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7924_), .Y(_7925_) );
	NAND3X1 NAND3X1_1712 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .B(_7923_), .C(_7925_), .Y(_7926_) );
	NAND3X1 NAND3X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7921_), .C(_7791_), .Y(_7927_) );
	INVX1 INVX1_1175 ( .gnd(gnd), .vdd(vdd), .A(_7924_), .Y(_7928_) );
	OAI21X1 OAI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7928_), .Y(_7930_) );
	NAND3X1 NAND3X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf2), .B(_7927_), .C(_7930_), .Y(_7931_) );
	NAND2X1 NAND2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_7926_), .B(_7931_), .Y(_7932_) );
	NAND3X1 NAND3X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_7917_), .B(_7920_), .C(_7932_), .Y(_7933_) );
	OAI21X1 OAI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf4), .B(_7450__bF_buf0), .C(_7345_), .Y(_7934_) );
	NAND2X1 NAND2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .B(_7346_), .Y(_7935_) );
	NAND2X1 NAND2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_7353_), .B(_7357_), .Y(_7936_) );
	INVX1 INVX1_1176 ( .gnd(gnd), .vdd(vdd), .A(_7936_), .Y(_7937_) );
	OAI21X1 OAI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_7937_), .B(_7476_), .C(_7441_), .Y(_7938_) );
	XNOR2X1 XNOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_7938_), .B(_7935_), .Y(_7939_) );
	NAND3X1 NAND3X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7939_), .C(_7791_), .Y(_7941_) );
	NAND3X1 NAND3X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf1), .B(_7941_), .C(_7934_), .Y(_7942_) );
	INVX1 INVX1_1177 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .Y(_7943_) );
	OAI21X1 OAI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf3), .B(_7450__bF_buf5), .C(_7943_), .Y(_7944_) );
	INVX1 INVX1_1178 ( .gnd(gnd), .vdd(vdd), .A(_7939_), .Y(_7945_) );
	NAND3X1 NAND3X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_7945_), .C(_7791_), .Y(_7946_) );
	NAND3X1 NAND3X1_1719 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .B(_7946_), .C(_7944_), .Y(_7947_) );
	XNOR2X1 XNOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_7306_), .B(_7937_), .Y(_7948_) );
	INVX1 INVX1_1179 ( .gnd(gnd), .vdd(vdd), .A(_7948_), .Y(_7949_) );
	NAND2X1 NAND2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_7949_), .B(divider_divuResult_5_bF_buf3), .Y(_7950_) );
	OAI21X1 OAI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_7355_), .B(divider_divuResult_6_bF_buf1), .C(_7350_), .Y(_7952_) );
	OAI21X1 OAI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf2), .B(_7450__bF_buf4), .C(_7952_), .Y(_7953_) );
	NAND3X1 NAND3X1_1720 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .B(_7953_), .C(_7950_), .Y(_7954_) );
	NAND2X1 NAND2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_7948_), .B(divider_divuResult_5_bF_buf2), .Y(_7955_) );
	INVX1 INVX1_1180 ( .gnd(gnd), .vdd(vdd), .A(_7952_), .Y(_7956_) );
	OAI21X1 OAI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf1), .B(_7450__bF_buf3), .C(_7956_), .Y(_7957_) );
	NAND3X1 NAND3X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_7957_), .C(_7955_), .Y(_7958_) );
	NAND2X1 NAND2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_7954_), .B(_7958_), .Y(_7959_) );
	NAND3X1 NAND3X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_7942_), .B(_7947_), .C(_7959_), .Y(_7960_) );
	NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_7933_), .B(_7960_), .Y(_7961_) );
	NAND3X1 NAND3X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_7909_), .B(_7961_), .C(_7840_), .Y(_7963_) );
	OAI21X1 OAI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_7943_), .B(divider_divuResult_5_bF_buf1), .C(_7941_), .Y(_7964_) );
	NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .B(_7964_), .Y(_7965_) );
	AOI21X1 AOI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(_7957_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .Y(_7966_) );
	OAI21X1 OAI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_7966_), .B(_7965_), .C(_7947_), .Y(_7967_) );
	INVX1 INVX1_1181 ( .gnd(gnd), .vdd(vdd), .A(_7917_), .Y(_7968_) );
	AOI21X1 AOI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_7930_), .B(_7927_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .Y(_7969_) );
	AOI21X1 AOI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .B(_7920_), .C(_7968_), .Y(_7970_) );
	OAI21X1 OAI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .B(_7933_), .C(_7970_), .Y(_7971_) );
	INVX1 INVX1_1182 ( .gnd(gnd), .vdd(vdd), .A(_7887_), .Y(_7972_) );
	AOI21X1 AOI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_7904_), .B(_7902_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .Y(_7974_) );
	OAI21X1 OAI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_7974_), .B(_7972_), .C(_7894_), .Y(_7975_) );
	OAI21X1 OAI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_7516_), .B(divider_divuResult_5_bF_buf0), .C(_7854_), .Y(_7976_) );
	INVX1 INVX1_1183 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .Y(_7977_) );
	OAI21X1 OAI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_7868_), .B(divider_divuResult_5_bF_buf6), .C(_7862_), .Y(_7978_) );
	OAI21X1 OAI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .B(_7978_), .C(_7855_), .Y(_7979_) );
	OAI21X1 OAI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf4), .B(_7977_), .C(_7979_), .Y(_7980_) );
	OAI21X1 OAI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_7872_), .B(_7975_), .C(_7980_), .Y(_7981_) );
	AOI21X1 AOI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_7971_), .B(_7909_), .C(_7981_), .Y(_7982_) );
	NAND2X1 NAND2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_7716_), .B(_7723_), .Y(_7983_) );
	AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .B(_7734_), .Y(_7985_) );
	NAND3X1 NAND3X1_1724 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .B(_7747_), .C(_7746_), .Y(_7986_) );
	AOI21X1 AOI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .B(_7744_), .C(_7508_), .Y(_7987_) );
	AOI21X1 AOI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_7163_), .B(_7165_), .C(divider_divuResult_5_bF_buf5), .Y(_7988_) );
	OAI21X1 OAI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_7988_), .B(_7987_), .C(_1494__bF_buf3), .Y(_7989_) );
	OAI21X1 OAI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_7740_), .B(_7751_), .C(divider_divuResult_5_bF_buf4), .Y(_7990_) );
	OAI21X1 OAI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf0), .B(_7450__bF_buf2), .C(_7750_), .Y(_7991_) );
	NAND3X1 NAND3X1_1725 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .B(_7991_), .C(_7990_), .Y(_7992_) );
	OAI21X1 OAI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_6315__bF_buf5), .B(_7450__bF_buf1), .C(_7749_), .Y(_7993_) );
	NAND3X1 NAND3X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf0), .B(_7993_), .C(_7754_), .Y(_7994_) );
	AOI22X1 AOI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(_7992_), .B(_7994_), .C(_7986_), .D(_7989_), .Y(_7996_) );
	NAND3X1 NAND3X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_7983_), .B(_7985_), .C(_7996_), .Y(_7997_) );
	INVX1 INVX1_1184 ( .gnd(gnd), .vdd(vdd), .A(_7997_), .Y(_7998_) );
	NAND3X1 NAND3X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_7672_), .B(_7699_), .C(_7998_), .Y(_7999_) );
	AOI21X1 AOI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7982_), .C(_7999_), .Y(_8000_) );
	OAI21X1 OAI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_7781_), .B(_8000_), .C(_7638_), .Y(_8001_) );
	AOI21X1 AOI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_8001_), .B(_7614_), .C(_2031_), .Y(divider_divuResult_4_) );
	AOI21X1 AOI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_7823_), .B(_7818_), .C(_2470__bF_buf3), .Y(_8002_) );
	OAI21X1 OAI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_7811_), .B(divider_divuResult_5_bF_buf3), .C(_7816_), .Y(_8003_) );
	NAND2X1 NAND2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf4), .B(_8003_), .Y(_8004_) );
	AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .B(_7817_), .Y(_8006_) );
	AOI21X1 AOI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_7797_), .B(_7796_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .Y(_8007_) );
	INVX1 INVX1_1185 ( .gnd(gnd), .vdd(vdd), .A(_7800_), .Y(_8008_) );
	AOI21X1 AOI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_7798_), .B(_8008_), .C(_8007_), .Y(_8009_) );
	OAI21X1 OAI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_8006_), .B(_8009_), .C(_8004_), .Y(_8010_) );
	INVX1 INVX1_1186 ( .gnd(gnd), .vdd(vdd), .A(_8010_), .Y(_8011_) );
	OAI21X1 OAI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_8002_), .B(_7834_), .C(_8011_), .Y(_8012_) );
	OAI21X1 OAI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7822_), .C(_7827_), .Y(_8013_) );
	NAND2X1 NAND2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_8013_), .Y(_8014_) );
	NAND3X1 NAND3X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_8014_), .C(_8010_), .Y(_8015_) );
	NAND2X1 NAND2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_8015_), .B(_8012_), .Y(_8017_) );
	NAND2X1 NAND2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_8017_), .B(divider_divuResult_4_bF_buf6), .Y(_8018_) );
	INVX8 INVX8_40 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .Y(_8019_) );
	INVX1 INVX1_1187 ( .gnd(gnd), .vdd(vdd), .A(_7627_), .Y(_8020_) );
	INVX1 INVX1_1188 ( .gnd(gnd), .vdd(vdd), .A(_7633_), .Y(_8021_) );
	OAI21X1 OAI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_8020_), .B(_8021_), .C(_7635_), .Y(_8022_) );
	NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_7579_), .B(_8022_), .Y(_8023_) );
	NAND2X1 NAND2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_7546_), .Y(_8024_) );
	NAND3X1 NAND3X1_1730 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf4), .B(_7660_), .C(_7658_), .Y(_8025_) );
	NAND2X1 NAND2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_7671_), .B(_7666_), .Y(_8026_) );
	NAND3X1 NAND3X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_8026_), .B(_7774_), .C(_8025_), .Y(_8028_) );
	AOI21X1 AOI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_7770_), .B(_7767_), .C(divider_absoluteValue_B_flipSign_result_17_bF_buf0), .Y(_8029_) );
	OAI22X1 OAI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_7694_), .B(_7696_), .C(_7685_), .D(_8029_), .Y(_8030_) );
	NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(_8028_), .Y(_8031_) );
	NAND2X1 NAND2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_7983_), .B(_7985_), .Y(_8032_) );
	INVX1 INVX1_1189 ( .gnd(gnd), .vdd(vdd), .A(_7758_), .Y(_8033_) );
	INVX1 INVX1_1190 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .Y(_8034_) );
	AOI21X1 AOI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_7983_), .B(_8034_), .C(_7760_), .Y(_8035_) );
	OAI21X1 OAI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_8032_), .B(_8033_), .C(_8035_), .Y(_8036_) );
	OAI21X1 OAI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_7673_), .B(divider_divuResult_5_bF_buf2), .C(_7770_), .Y(_8037_) );
	NAND2X1 NAND2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .B(_8037_), .Y(_8039_) );
	INVX1 INVX1_1191 ( .gnd(gnd), .vdd(vdd), .A(_7772_), .Y(_8040_) );
	OAI21X1 OAI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_7765_), .B(_8040_), .C(_8039_), .Y(_8041_) );
	AOI21X1 AOI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_7658_), .B(_7660_), .C(divider_absoluteValue_B_flipSign_result_19_bF_buf3), .Y(_8042_) );
	NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf4), .B(_7777_), .Y(_8043_) );
	AOI21X1 AOI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_8025_), .B(_8043_), .C(_8042_), .Y(_8044_) );
	OAI21X1 OAI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_8041_), .B(_8028_), .C(_8044_), .Y(_8045_) );
	AOI21X1 AOI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_8031_), .B(_8036_), .C(_8045_), .Y(_8046_) );
	OAI21X1 OAI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_8024_), .B(_8046_), .C(_7614_), .Y(_8047_) );
	NOR3X1 NOR3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_8030_), .B(_7997_), .C(_8028_), .Y(_8048_) );
	NAND3X1 NAND3X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_7546_), .C(_8048_), .Y(_8050_) );
	AOI21X1 AOI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7982_), .C(_8050_), .Y(_8051_) );
	OAI21X1 OAI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .B(_8047_), .C(_8019__bF_buf3), .Y(_8052_) );
	NAND3X1 NAND3X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_7826_), .B(_7827_), .C(_8052__bF_buf6), .Y(_8053_) );
	NAND3X1 NAND3X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_8053_), .C(_8018_), .Y(_8054_) );
	INVX1 INVX1_1192 ( .gnd(gnd), .vdd(vdd), .A(_8054_), .Y(_8055_) );
	INVX1 INVX1_1193 ( .gnd(gnd), .vdd(vdd), .A(_8017_), .Y(_8056_) );
	NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_8056_), .B(_8052__bF_buf5), .Y(_8057_) );
	NAND2X1 NAND2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_7781_), .B(_7638_), .Y(_8058_) );
	NAND2X1 NAND2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_7982_), .B(_7963_), .Y(_8059_) );
	NAND3X1 NAND3X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .B(_8059_), .C(_7638_), .Y(_8061_) );
	NAND3X1 NAND3X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_7614_), .B(_8058_), .C(_8061_), .Y(_8062_) );
	AOI21X1 AOI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_8062__bF_buf3), .B(_8019__bF_buf2), .C(_8013_), .Y(_8063_) );
	OAI21X1 OAI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .B(_8057_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf5), .Y(_8064_) );
	XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_8009_), .B(_8006_), .Y(_8065_) );
	INVX1 INVX1_1194 ( .gnd(gnd), .vdd(vdd), .A(_8065_), .Y(_8066_) );
	NAND3X1 NAND3X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf1), .B(_8066_), .C(_8062__bF_buf2), .Y(_8067_) );
	OAI21X1 OAI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_8003_), .B(divider_divuResult_4_bF_buf5), .C(_8067_), .Y(_8068_) );
	NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf0), .B(_8068_), .Y(_8069_) );
	AOI21X1 AOI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_8069_), .B(_8064_), .C(_8055_), .Y(_8070_) );
	NAND3X1 NAND3X1_1738 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf4), .B(_8053_), .C(_8018_), .Y(_8072_) );
	OAI21X1 OAI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .B(_8057_), .C(_1735__bF_buf0), .Y(_8073_) );
	INVX1 INVX1_1195 ( .gnd(gnd), .vdd(vdd), .A(_8003_), .Y(_8074_) );
	NAND2X1 NAND2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_8074_), .B(_8052__bF_buf4), .Y(_8075_) );
	NAND3X1 NAND3X1_1739 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf7), .B(_8067_), .C(_8075_), .Y(_8076_) );
	NAND3X1 NAND3X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf0), .B(_8065_), .C(_8062__bF_buf1), .Y(_8077_) );
	NAND2X1 NAND2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_8003_), .B(_8052__bF_buf3), .Y(_8078_) );
	NAND3X1 NAND3X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_8077_), .C(_8078_), .Y(_8079_) );
	AOI22X1 AOI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(_8076_), .B(_8079_), .C(_8072_), .D(_8073_), .Y(_8080_) );
	XNOR2X1 XNOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_7799_), .B(_7800_), .Y(_8081_) );
	INVX1 INVX1_1196 ( .gnd(gnd), .vdd(vdd), .A(_8081_), .Y(_8083_) );
	NAND3X1 NAND3X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf3), .B(_8083_), .C(_8062__bF_buf0), .Y(_8084_) );
	OAI21X1 OAI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_5_), .B(divider_divuResult_5_bF_buf1), .C(_7792_), .Y(_8085_) );
	NAND2X1 NAND2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_8085_), .B(_8052__bF_buf2), .Y(_8086_) );
	AOI21X1 AOI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_8086_), .B(_8084_), .C(_2547__bF_buf3), .Y(_8087_) );
	NAND3X1 NAND3X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf2), .B(_7803_), .C(_8062__bF_buf3), .Y(_8088_) );
	NAND2X1 NAND2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_7801_), .B(_8052__bF_buf1), .Y(_8089_) );
	NAND3X1 NAND3X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf1), .B(_8088_), .C(_8089_), .Y(_8090_) );
	NAND3X1 NAND3X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf1), .B(_8081_), .C(_8062__bF_buf2), .Y(_8091_) );
	OAI21X1 OAI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_8085_), .B(divider_divuResult_4_bF_buf4), .C(_8091_), .Y(_8092_) );
	NAND2X1 NAND2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf2), .B(_8092_), .Y(_8094_) );
	OAI21X1 OAI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_8087_), .B(_8090_), .C(_8094_), .Y(_8095_) );
	NAND2X1 NAND2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_8095_), .B(_8080_), .Y(_8096_) );
	NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_3_), .B(_1746__bF_buf5), .Y(_8097_) );
	INVX1 INVX1_1197 ( .gnd(gnd), .vdd(vdd), .A(_8097_), .Y(_8098_) );
	NAND3X1 NAND3X1_1746 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .B(_8088_), .C(_8089_), .Y(_8099_) );
	NAND2X1 NAND2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf4), .B(_8019__bF_buf0), .Y(_8100_) );
	INVX1 INVX1_1198 ( .gnd(gnd), .vdd(vdd), .A(_8100_), .Y(_8101_) );
	OAI21X1 OAI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .B(_8047_), .C(_8101_), .Y(_8102_) );
	NAND2X1 NAND2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_4_), .B(_8102_), .Y(_8103_) );
	NAND3X1 NAND3X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_7801_), .B(_8101_), .C(_8062__bF_buf1), .Y(_8105_) );
	NAND3X1 NAND3X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf0), .B(_8105_), .C(_8103_), .Y(_8106_) );
	NAND3X1 NAND3X1_1749 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf7), .B(_8084_), .C(_8086_), .Y(_8107_) );
	INVX1 INVX1_1199 ( .gnd(gnd), .vdd(vdd), .A(_8085_), .Y(_8108_) );
	NAND2X1 NAND2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_8108_), .B(_8052__bF_buf0), .Y(_8109_) );
	NAND3X1 NAND3X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf1), .B(_8091_), .C(_8109_), .Y(_8110_) );
	AOI22X1 AOI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(_8099_), .B(_8106_), .C(_8107_), .D(_8110_), .Y(_8111_) );
	NAND3X1 NAND3X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_8111_), .C(_8080_), .Y(_8112_) );
	NAND3X1 NAND3X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_8070_), .B(_8096_), .C(_8112_), .Y(_8113_) );
	NAND2X1 NAND2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_7855_), .B(_7860_), .Y(_8114_) );
	INVX1 INVX1_1200 ( .gnd(gnd), .vdd(vdd), .A(_8114_), .Y(_8116_) );
	NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .B(_7978_), .Y(_8117_) );
	INVX1 INVX1_1201 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .Y(_8118_) );
	NAND2X1 NAND2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_7887_), .B(_7894_), .Y(_8119_) );
	INVX1 INVX1_1202 ( .gnd(gnd), .vdd(vdd), .A(_7974_), .Y(_8120_) );
	OAI21X1 OAI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_8119_), .B(_8120_), .C(_7887_), .Y(_8121_) );
	NAND2X1 NAND2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_7917_), .B(_7920_), .Y(_8122_) );
	AOI21X1 AOI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_7926_), .B(_7931_), .C(_8122_), .Y(_8123_) );
	NAND2X1 NAND2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_7942_), .B(_7947_), .Y(_8124_) );
	OAI21X1 OAI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7949_), .C(_7957_), .Y(_8125_) );
	NAND2X1 NAND2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf7), .B(_8125_), .Y(_8127_) );
	OAI21X1 OAI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_8127_), .B(_8124_), .C(_7942_), .Y(_8128_) );
	INVX1 INVX1_1203 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .Y(_8129_) );
	OAI21X1 OAI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_8129_), .B(_8122_), .C(_7917_), .Y(_8130_) );
	AOI21X1 AOI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_8123_), .B(_8128_), .C(_8130_), .Y(_8131_) );
	NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_7833_), .B(_7834_), .Y(_8132_) );
	OAI21X1 OAI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_8006_), .B(_8009_), .C(_8132_), .Y(_8133_) );
	NAND3X1 NAND3X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_8133_), .C(_7961_), .Y(_8134_) );
	AOI21X1 AOI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_8134_), .B(_8131_), .C(_7908_), .Y(_8135_) );
	OAI21X1 OAI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_8121_), .B(_8135_), .C(_7871_), .Y(_8136_) );
	NAND3X1 NAND3X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_8116_), .B(_8118_), .C(_8136_), .Y(_8138_) );
	AOI21X1 AOI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .B(_7905_), .C(_8119_), .Y(_8139_) );
	OAI21X1 OAI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_8004_), .B(_8002_), .C(_8014_), .Y(_8140_) );
	AOI21X1 AOI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_7838_), .B(_7829_), .C(_8140_), .Y(_8141_) );
	AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_7920_), .B(_7917_), .Y(_8142_) );
	AOI21X1 AOI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_7954_), .B(_7958_), .C(_8124_), .Y(_8143_) );
	NAND3X1 NAND3X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_8142_), .B(_7932_), .C(_8143_), .Y(_8144_) );
	AOI21X1 AOI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_7831_), .B(_8141_), .C(_8144_), .Y(_8145_) );
	OAI21X1 OAI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_7971_), .B(_8145_), .C(_8139_), .Y(_8146_) );
	AOI22X1 AOI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(_7865_), .B(_7870_), .C(_7975_), .D(_8146_), .Y(_8147_) );
	OAI21X1 OAI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .B(_8147_), .C(_8114_), .Y(_8149_) );
	AOI21X1 AOI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_8149_), .B(_8138_), .C(_8052__bF_buf6), .Y(_8150_) );
	AOI21X1 AOI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_8062__bF_buf0), .B(_8019__bF_buf3), .C(_7976_), .Y(_8151_) );
	OAI21X1 OAI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_8151_), .B(_8150_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .Y(_8152_) );
	AOI21X1 AOI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_8062__bF_buf3), .B(_8019__bF_buf2), .C(_7977_), .Y(_8153_) );
	OAI21X1 OAI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .B(_8147_), .C(_8116_), .Y(_8154_) );
	NAND3X1 NAND3X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_8114_), .B(_8118_), .C(_8136_), .Y(_8155_) );
	AOI21X1 AOI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_8154_), .B(_8155_), .C(_8052__bF_buf5), .Y(_8156_) );
	OAI21X1 OAI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_8153_), .B(_8156_), .C(_1484__bF_buf4), .Y(_8157_) );
	INVX1 INVX1_1204 ( .gnd(gnd), .vdd(vdd), .A(_7871_), .Y(_8158_) );
	NAND3X1 NAND3X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_8158_), .B(_7975_), .C(_8146_), .Y(_8160_) );
	NAND2X1 NAND2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_8160_), .B(_8136_), .Y(_8161_) );
	NAND3X1 NAND3X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf1), .B(_8161_), .C(_8062__bF_buf2), .Y(_8162_) );
	NAND2X1 NAND2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_7978_), .B(_8052__bF_buf4), .Y(_8163_) );
	NAND3X1 NAND3X1_1759 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .B(_8162_), .C(_8163_), .Y(_8164_) );
	AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_8136_), .B(_8160_), .Y(_8165_) );
	NAND3X1 NAND3X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf0), .B(_8062__bF_buf1), .C(_8165_), .Y(_8166_) );
	INVX1 INVX1_1205 ( .gnd(gnd), .vdd(vdd), .A(_7978_), .Y(_8167_) );
	NAND2X1 NAND2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_8167_), .B(_8052__bF_buf3), .Y(_8168_) );
	NAND3X1 NAND3X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf3), .B(_8168_), .C(_8166_), .Y(_8169_) );
	AOI22X1 AOI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(_8164_), .B(_8169_), .C(_8152_), .D(_8157_), .Y(_8171_) );
	NAND3X1 NAND3X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_7889_), .B(_7893_), .C(_8052__bF_buf2), .Y(_8172_) );
	INVX1 INVX1_1206 ( .gnd(gnd), .vdd(vdd), .A(_8119_), .Y(_8173_) );
	AOI22X1 AOI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .B(_7905_), .C(_8131_), .D(_8134_), .Y(_8174_) );
	OAI21X1 OAI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_7974_), .B(_8174_), .C(_8173_), .Y(_8175_) );
	OAI21X1 OAI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_7971_), .B(_8145_), .C(_7906_), .Y(_8176_) );
	NAND3X1 NAND3X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_8119_), .B(_8120_), .C(_8176_), .Y(_8177_) );
	NAND2X1 NAND2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_8177_), .B(_8175_), .Y(_8178_) );
	NAND3X1 NAND3X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf3), .B(_8178_), .C(_8062__bF_buf0), .Y(_8179_) );
	NAND3X1 NAND3X1_1765 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .B(_8179_), .C(_8172_), .Y(_8180_) );
	OAI21X1 OAI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7884_), .C(_7889_), .Y(_8182_) );
	NAND2X1 NAND2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_8182_), .B(_8052__bF_buf1), .Y(_8183_) );
	AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_8175_), .B(_8177_), .Y(_8184_) );
	NAND2X1 NAND2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_8184_), .B(divider_divuResult_4_bF_buf3), .Y(_8185_) );
	NAND3X1 NAND3X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf1), .B(_8183_), .C(_8185_), .Y(_8186_) );
	NAND2X1 NAND2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_8133_), .Y(_8187_) );
	OAI21X1 OAI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_8144_), .B(_8187_), .C(_8131_), .Y(_8188_) );
	NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_7906_), .B(_8188_), .Y(_8189_) );
	NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_8174_), .B(_8189_), .Y(_8190_) );
	INVX1 INVX1_1207 ( .gnd(gnd), .vdd(vdd), .A(_8190_), .Y(_8191_) );
	NAND3X1 NAND3X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf2), .B(_8191_), .C(_8062__bF_buf3), .Y(_8193_) );
	NAND3X1 NAND3X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_7902_), .B(_7904_), .C(_8052__bF_buf0), .Y(_8194_) );
	NAND3X1 NAND3X1_1769 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_8193_), .C(_8194_), .Y(_8195_) );
	NAND3X1 NAND3X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf1), .B(_8190_), .C(_8062__bF_buf2), .Y(_8196_) );
	OAI21X1 OAI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .B(_7897_), .C(_7902_), .Y(_8197_) );
	NAND2X1 NAND2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_8197_), .B(_8052__bF_buf6), .Y(_8198_) );
	NAND3X1 NAND3X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf0), .B(_8196_), .C(_8198_), .Y(_8199_) );
	AOI22X1 AOI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(_8195_), .B(_8199_), .C(_8180_), .D(_8186_), .Y(_8200_) );
	NAND2X1 NAND2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_8200_), .B(_8171_), .Y(_8201_) );
	NAND2X1 NAND2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_7919_), .B(_8052__bF_buf5), .Y(_8202_) );
	OAI21X1 OAI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .B(_8187_), .C(_7967_), .Y(_8204_) );
	AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_8204_), .B(_7932_), .Y(_8205_) );
	OAI21X1 OAI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .B(_8205_), .C(_8142_), .Y(_8206_) );
	NAND2X1 NAND2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_7932_), .B(_8204_), .Y(_8207_) );
	NAND3X1 NAND3X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_8122_), .B(_8129_), .C(_8207_), .Y(_8208_) );
	NAND2X1 NAND2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_8208_), .B(_8206_), .Y(_8209_) );
	NAND3X1 NAND3X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf0), .B(_8062__bF_buf1), .C(_8209_), .Y(_8210_) );
	NAND3X1 NAND3X1_1774 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .B(_8202_), .C(_8210_), .Y(_8211_) );
	AOI22X1 AOI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(_7910_), .B(_7916_), .C(_8019__bF_buf3), .D(_8062__bF_buf0), .Y(_8212_) );
	AOI21X1 AOI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_8206_), .B(_8208_), .C(_8052__bF_buf4), .Y(_8213_) );
	OAI21X1 OAI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_8212_), .B(_8213_), .C(_7204__bF_buf0), .Y(_8215_) );
	NAND2X1 NAND2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_8211_), .B(_8215_), .Y(_8216_) );
	XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_8204_), .B(_7932_), .Y(_8217_) );
	INVX1 INVX1_1208 ( .gnd(gnd), .vdd(vdd), .A(_8217_), .Y(_8218_) );
	NAND3X1 NAND3X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf2), .B(_8218_), .C(_8062__bF_buf3), .Y(_8219_) );
	OAI21X1 OAI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_7924_), .B(divider_divuResult_5_bF_buf0), .C(_7927_), .Y(_8220_) );
	INVX1 INVX1_1209 ( .gnd(gnd), .vdd(vdd), .A(_8220_), .Y(_8221_) );
	NAND2X1 NAND2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_8221_), .B(_8052__bF_buf3), .Y(_8222_) );
	NAND3X1 NAND3X1_1776 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .B(_8219_), .C(_8222_), .Y(_8223_) );
	NAND3X1 NAND3X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf1), .B(_8217_), .C(_8062__bF_buf2), .Y(_8224_) );
	NAND2X1 NAND2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_8220_), .B(_8052__bF_buf2), .Y(_8226_) );
	NAND3X1 NAND3X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf5), .B(_8224_), .C(_8226_), .Y(_8227_) );
	NAND2X1 NAND2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_8223_), .B(_8227_), .Y(_8228_) );
	NAND2X1 NAND2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_7964_), .B(_8052__bF_buf1), .Y(_8229_) );
	INVX1 INVX1_1210 ( .gnd(gnd), .vdd(vdd), .A(_7959_), .Y(_8230_) );
	OAI21X1 OAI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_8230_), .B(_8187_), .C(_8127_), .Y(_8231_) );
	NAND3X1 NAND3X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_7942_), .B(_7947_), .C(_8231_), .Y(_8232_) );
	INVX1 INVX1_1211 ( .gnd(gnd), .vdd(vdd), .A(_8231_), .Y(_8233_) );
	NAND2X1 NAND2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_8124_), .B(_8233_), .Y(_8234_) );
	NAND2X1 NAND2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_8232_), .B(_8234_), .Y(_8235_) );
	NAND3X1 NAND3X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf0), .B(_8235_), .C(_8062__bF_buf1), .Y(_8237_) );
	NAND3X1 NAND3X1_1781 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_8237_), .C(_8229_), .Y(_8238_) );
	INVX1 INVX1_1212 ( .gnd(gnd), .vdd(vdd), .A(_7964_), .Y(_8239_) );
	NAND2X1 NAND2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_8239_), .B(_8052__bF_buf0), .Y(_8240_) );
	AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_8234_), .B(_8232_), .Y(_8241_) );
	NAND3X1 NAND3X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf3), .B(_8241_), .C(_8062__bF_buf0), .Y(_8242_) );
	NAND3X1 NAND3X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_8242_), .C(_8240_), .Y(_8243_) );
	XNOR2X1 XNOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_8187_), .B(_7959_), .Y(_8244_) );
	INVX1 INVX1_1213 ( .gnd(gnd), .vdd(vdd), .A(_8244_), .Y(_8245_) );
	NAND3X1 NAND3X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf2), .B(_8245_), .C(_8062__bF_buf3), .Y(_8246_) );
	NAND3X1 NAND3X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(_7957_), .C(_8052__bF_buf6), .Y(_8248_) );
	NAND3X1 NAND3X1_1786 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf7), .B(_8246_), .C(_8248_), .Y(_8249_) );
	NAND3X1 NAND3X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_8019__bF_buf1), .B(_8244_), .C(_8062__bF_buf2), .Y(_8250_) );
	NAND2X1 NAND2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .B(_8052__bF_buf5), .Y(_8251_) );
	NAND3X1 NAND3X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf0), .B(_8250_), .C(_8251_), .Y(_8252_) );
	AOI22X1 AOI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(_8238_), .B(_8243_), .C(_8249_), .D(_8252_), .Y(_8253_) );
	NAND3X1 NAND3X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_8228_), .B(_8216_), .C(_8253_), .Y(_8254_) );
	NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_8254_), .B(_8201_), .Y(_8255_) );
	OAI21X1 OAI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_8153_), .B(_8156_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .Y(_8256_) );
	NAND2X1 NAND2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_8138_), .B(_8149_), .Y(_8257_) );
	NAND2X1 NAND2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .B(_8052__bF_buf4), .Y(_8259_) );
	OAI21X1 OAI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_8052__bF_buf3), .B(_8257_), .C(_8259_), .Y(_8260_) );
	OAI21X1 OAI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_8052__bF_buf2), .B(_8161_), .C(_8168_), .Y(_8261_) );
	NAND2X1 NAND2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf2), .B(_8261_), .Y(_8262_) );
	OAI21X1 OAI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .B(_8260_), .C(_8262_), .Y(_8263_) );
	AOI21X1 AOI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_8172_), .B(_8179_), .C(_10678__bF_buf0), .Y(_8264_) );
	NAND3X1 NAND3X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf5), .B(_8179_), .C(_8172_), .Y(_8265_) );
	NAND3X1 NAND3X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf6), .B(_8193_), .C(_8194_), .Y(_8266_) );
	AOI21X1 AOI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .B(_8265_), .C(_8264_), .Y(_8267_) );
	AOI22X1 AOI22X1_179 ( .gnd(gnd), .vdd(vdd), .A(_8171_), .B(_8267_), .C(_8256_), .D(_8263_), .Y(_8268_) );
	OAI21X1 OAI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_8212_), .B(_8213_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .Y(_8270_) );
	AOI22X1 AOI22X1_180 ( .gnd(gnd), .vdd(vdd), .A(_8223_), .B(_8227_), .C(_8211_), .D(_8215_), .Y(_8271_) );
	NAND3X1 NAND3X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf5), .B(_8202_), .C(_8210_), .Y(_8272_) );
	OAI21X1 OAI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_8220_), .B(divider_divuResult_4_bF_buf2), .C(_8219_), .Y(_8273_) );
	OAI21X1 OAI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_8273_), .C(_8272_), .Y(_8274_) );
	NAND3X1 NAND3X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf0), .B(_8237_), .C(_8229_), .Y(_8275_) );
	AOI21X1 AOI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_8229_), .B(_8237_), .C(_4999__bF_buf6), .Y(_8276_) );
	NAND3X1 NAND3X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf7), .B(_8246_), .C(_8248_), .Y(_8277_) );
	AOI21X1 AOI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_8277_), .B(_8275_), .C(_8276_), .Y(_8278_) );
	AOI22X1 AOI22X1_181 ( .gnd(gnd), .vdd(vdd), .A(_8270_), .B(_8274_), .C(_8278_), .D(_8271_), .Y(_8279_) );
	OAI21X1 OAI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_8201_), .B(_8279_), .C(_8268_), .Y(_8281_) );
	AOI21X1 AOI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_8113_), .B(_8255_), .C(_8281_), .Y(_8282_) );
	OAI21X1 OAI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_7451_), .B(divider_divuResult_4_bF_buf1), .C(_2229__bF_buf0), .Y(_8283_) );
	NAND2X1 NAND2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .B(_8283_), .Y(_8284_) );
	OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_8283_), .B(divider_absoluteValue_B_flipSign_result_28_), .Y(_8285_) );
	NAND2X1 NAND2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_8284_), .B(_8285_), .Y(_8286_) );
	AOI21X1 AOI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_7865_), .B(_7870_), .C(_8114_), .Y(_8287_) );
	NAND2X1 NAND2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_8139_), .B(_8287_), .Y(_8288_) );
	NOR3X1 NOR3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_8288_), .B(_8144_), .C(_8187_), .Y(_8289_) );
	AOI22X1 AOI22X1_182 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_7860_), .C(_8287_), .D(_8121_), .Y(_8290_) );
	OAI21X1 OAI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_8288_), .B(_8131_), .C(_8290_), .Y(_8292_) );
	OAI21X1 OAI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_8292_), .B(_8289_), .C(_8048_), .Y(_8293_) );
	AOI21X1 AOI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_8293_), .B(_8046_), .C(_7637_), .Y(_8294_) );
	OAI21X1 OAI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_7606_), .B(_8294_), .C(_7623_), .Y(_8295_) );
	AOI22X1 AOI22X1_183 ( .gnd(gnd), .vdd(vdd), .A(_7616_), .B(_7617_), .C(_7609_), .D(_8295_), .Y(_8296_) );
	NAND2X1 NAND2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_7617_), .B(_7616_), .Y(_8297_) );
	INVX1 INVX1_1214 ( .gnd(gnd), .vdd(vdd), .A(_7609_), .Y(_8298_) );
	INVX1 INVX1_1215 ( .gnd(gnd), .vdd(vdd), .A(_7606_), .Y(_8299_) );
	OAI21X1 OAI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_7781_), .B(_8000_), .C(_8023_), .Y(_8300_) );
	AOI21X1 AOI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_8300_), .B(_8299_), .C(_7545_), .Y(_8301_) );
	NOR3X1 NOR3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_8297_), .B(_8298_), .C(_8301_), .Y(_8303_) );
	OAI21X1 OAI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_8303_), .B(_8296_), .C(divider_divuResult_4_bF_buf0), .Y(_8304_) );
	NAND2X1 NAND2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_7502_), .B(_7501_), .Y(_8305_) );
	OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf6), .B(_8305_), .Y(_8306_) );
	NAND3X1 NAND3X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_8306_), .C(_8304_), .Y(_8307_) );
	OAI21X1 OAI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_8298_), .B(_8301_), .C(_8297_), .Y(_8308_) );
	INVX1 INVX1_1216 ( .gnd(gnd), .vdd(vdd), .A(_8297_), .Y(_8309_) );
	NAND3X1 NAND3X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_8309_), .B(_7609_), .C(_8295_), .Y(_8310_) );
	NAND3X1 NAND3X1_1797 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf5), .B(_8308_), .C(_8310_), .Y(_8311_) );
	NAND2X1 NAND2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_8305_), .B(_8052__bF_buf1), .Y(_8312_) );
	NAND3X1 NAND3X1_1798 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_8312_), .C(_8311_), .Y(_8314_) );
	NAND3X1 NAND3X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_8286_), .B(_8314_), .C(_8307_), .Y(_8315_) );
	OAI21X1 OAI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_7528_), .B(_7531_), .C(_8052__bF_buf0), .Y(_8316_) );
	NAND2X1 NAND2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_7619_), .B(_7620_), .Y(_8317_) );
	OAI21X1 OAI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_7606_), .B(_8294_), .C(_7543_), .Y(_8318_) );
	NAND3X1 NAND3X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .B(_7537_), .C(_8318_), .Y(_8319_) );
	INVX1 INVX1_1217 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .Y(_8320_) );
	AOI21X1 AOI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_8300_), .B(_8299_), .C(_7622_), .Y(_8321_) );
	OAI21X1 OAI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_7608_), .B(_8321_), .C(_8320_), .Y(_8322_) );
	NAND3X1 NAND3X1_1801 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf4), .B(_8322_), .C(_8319_), .Y(_8323_) );
	NAND3X1 NAND3X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_8316_), .C(_8323_), .Y(_8325_) );
	INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(_8316_), .Y(_8326_) );
	OAI21X1 OAI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_7608_), .B(_8321_), .C(_8317_), .Y(_8327_) );
	NAND3X1 NAND3X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_8320_), .B(_7537_), .C(_8318_), .Y(_8328_) );
	AOI21X1 AOI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .B(_8327_), .C(_8052__bF_buf6), .Y(_8329_) );
	OAI21X1 OAI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_8326_), .B(_8329_), .C(divider_absoluteValue_B_flipSign_result_26_bF_buf2), .Y(_8330_) );
	NAND3X1 NAND3X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_7622_), .B(_8299_), .C(_8300_), .Y(_8331_) );
	INVX1 INVX1_1218 ( .gnd(gnd), .vdd(vdd), .A(_8331_), .Y(_8332_) );
	OAI21X1 OAI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_8321_), .B(_8332_), .C(divider_divuResult_4_bF_buf3), .Y(_8333_) );
	OAI21X1 OAI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_7461_), .B(divider_divuResult_5_bF_buf6), .C(_7540_), .Y(_8334_) );
	OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf2), .B(_8334_), .Y(_8335_) );
	NAND3X1 NAND3X1_1805 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_8335_), .C(_8333_), .Y(_8336_) );
	NAND3X1 NAND3X1_1806 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf1), .B(_8331_), .C(_8318_), .Y(_8337_) );
	NAND2X1 NAND2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_8334_), .B(_8052__bF_buf5), .Y(_8338_) );
	NAND3X1 NAND3X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_8338_), .C(_8337_), .Y(_8339_) );
	NAND2X1 NAND2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_8339_), .B(_8336_), .Y(_8340_) );
	NAND3X1 NAND3X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_8325_), .B(_8340_), .C(_8330_), .Y(_8341_) );
	NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8341_), .Y(_8342_) );
	OAI21X1 OAI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_7560_), .B(divider_divuResult_5_bF_buf5), .C(_7558_), .Y(_8343_) );
	NAND2X1 NAND2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_8343_), .B(_8052__bF_buf4), .Y(_8344_) );
	INVX1 INVX1_1219 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .Y(_8347_) );
	INVX1 INVX1_1220 ( .gnd(gnd), .vdd(vdd), .A(_7601_), .Y(_8348_) );
	AOI21X1 AOI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_8293_), .B(_8046_), .C(_8022_), .Y(_8349_) );
	OAI21X1 OAI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_8348_), .B(_8349_), .C(_7578_), .Y(_8350_) );
	NAND3X1 NAND3X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_7625_), .B(_8347_), .C(_8350_), .Y(_8351_) );
	INVX1 INVX1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7625_), .Y(_8352_) );
	INVX1 INVX1_1222 ( .gnd(gnd), .vdd(vdd), .A(_7578_), .Y(_8353_) );
	OAI21X1 OAI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_7781_), .B(_8000_), .C(_7636_), .Y(_8354_) );
	AOI21X1 AOI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_8354_), .B(_7601_), .C(_8353_), .Y(_8355_) );
	OAI21X1 OAI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .B(_8355_), .C(_8352_), .Y(_8356_) );
	NAND3X1 NAND3X1_1810 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf0), .B(_8356_), .C(_8351_), .Y(_8358_) );
	NAND3X1 NAND3X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf3), .B(_8344_), .C(_8358_), .Y(_8359_) );
	OAI21X1 OAI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_7604_), .B(_8355_), .C(_7625_), .Y(_8360_) );
	NAND3X1 NAND3X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_8352_), .B(_8347_), .C(_8350_), .Y(_8361_) );
	NAND3X1 NAND3X1_1813 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf6), .B(_8360_), .C(_8361_), .Y(_8362_) );
	INVX1 INVX1_1223 ( .gnd(gnd), .vdd(vdd), .A(_8343_), .Y(_8363_) );
	NAND2X1 NAND2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_8363_), .B(_8052__bF_buf3), .Y(_8364_) );
	NAND3X1 NAND3X1_1814 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf1), .B(_8364_), .C(_8362_), .Y(_8365_) );
	NAND3X1 NAND3X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_8353_), .B(_7601_), .C(_8354_), .Y(_8366_) );
	INVX1 INVX1_1224 ( .gnd(gnd), .vdd(vdd), .A(_8366_), .Y(_8367_) );
	OAI21X1 OAI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_8355_), .B(_8367_), .C(divider_divuResult_4_bF_buf5), .Y(_8369_) );
	OAI21X1 OAI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_7573_), .B(_7575_), .C(_8052__bF_buf2), .Y(_8370_) );
	NAND3X1 NAND3X1_1816 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf1), .B(_8370_), .C(_8369_), .Y(_8371_) );
	AOI21X1 AOI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_8350_), .B(_8366_), .C(_8052__bF_buf1), .Y(_8372_) );
	INVX1 INVX1_1225 ( .gnd(gnd), .vdd(vdd), .A(_7603_), .Y(_8373_) );
	NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .B(divider_divuResult_4_bF_buf4), .Y(_8374_) );
	OAI21X1 OAI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_8374_), .B(_8372_), .C(_5516__bF_buf1), .Y(_8375_) );
	NAND2X1 NAND2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_8371_), .B(_8375_), .Y(_8376_) );
	NAND3X1 NAND3X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_8359_), .B(_8365_), .C(_8376_), .Y(_8377_) );
	OAI21X1 OAI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_7781_), .B(_8000_), .C(_7635_), .Y(_8378_) );
	INVX1 INVX1_1226 ( .gnd(gnd), .vdd(vdd), .A(_8378_), .Y(_8380_) );
	NAND2X1 NAND2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_8046_), .B(_8293_), .Y(_8381_) );
	NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_7635_), .B(_8381_), .Y(_8382_) );
	OAI21X1 OAI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_8380_), .B(_8382_), .C(divider_divuResult_4_bF_buf3), .Y(_8383_) );
	OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf2), .B(_7597_), .Y(_8384_) );
	NAND3X1 NAND3X1_1818 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf1), .B(_8383_), .C(_8384_), .Y(_8385_) );
	OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_8381_), .B(_7635_), .Y(_8386_) );
	AOI21X1 AOI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_8386_), .B(_8378_), .C(_8052__bF_buf0), .Y(_8387_) );
	NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_7597_), .B(divider_divuResult_4_bF_buf1), .Y(_8388_) );
	OAI21X1 OAI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_8388_), .B(_8387_), .C(_4424__bF_buf1), .Y(_8389_) );
	NAND2X1 NAND2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_8385_), .B(_8389_), .Y(_8391_) );
	NAND2X1 NAND2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_7592_), .B(_8052__bF_buf6), .Y(_8392_) );
	NAND3X1 NAND3X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_7634_), .C(_8378_), .Y(_8393_) );
	INVX1 INVX1_1227 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .Y(_8394_) );
	NAND2X1 NAND2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_8378_), .Y(_8395_) );
	NAND2X1 NAND2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_8394_), .B(_8395_), .Y(_8396_) );
	NAND3X1 NAND3X1_1820 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf0), .B(_8393_), .C(_8396_), .Y(_8397_) );
	NAND3X1 NAND3X1_1821 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf0), .B(_8392_), .C(_8397_), .Y(_8398_) );
	INVX1 INVX1_1228 ( .gnd(gnd), .vdd(vdd), .A(_8392_), .Y(_8399_) );
	OAI21X1 OAI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_8020_), .B(_8021_), .C(_8395_), .Y(_8400_) );
	NAND3X1 NAND3X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_8394_), .C(_8378_), .Y(_8402_) );
	AOI21X1 AOI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_8400_), .B(_8402_), .C(_8052__bF_buf5), .Y(_8403_) );
	OAI21X1 OAI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_8399_), .B(_8403_), .C(_4881__bF_buf1), .Y(_8404_) );
	NAND2X1 NAND2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_8398_), .B(_8404_), .Y(_8405_) );
	NAND2X1 NAND2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_8391_), .B(_8405_), .Y(_8406_) );
	NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_8377_), .B(_8406_), .Y(_8407_) );
	OAI21X1 OAI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_7659_), .B(divider_divuResult_5_bF_buf4), .C(_7653_), .Y(_8408_) );
	NAND2X1 NAND2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_8408_), .B(_8052__bF_buf4), .Y(_8409_) );
	NAND2X1 NAND2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .B(_7661_), .Y(_8410_) );
	OAI21X1 OAI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_8292_), .B(_8289_), .C(_7998_), .Y(_8411_) );
	AOI21X1 AOI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_8411_), .B(_7763_), .C(_8030_), .Y(_8413_) );
	OAI21X1 OAI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_7773_), .B(_8413_), .C(_8026_), .Y(_8414_) );
	NAND3X1 NAND3X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_8410_), .B(_7778_), .C(_8414_), .Y(_8415_) );
	INVX1 INVX1_1229 ( .gnd(gnd), .vdd(vdd), .A(_8410_), .Y(_8416_) );
	INVX1 INVX1_1230 ( .gnd(gnd), .vdd(vdd), .A(_8026_), .Y(_8417_) );
	AOI21X1 AOI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7982_), .C(_7997_), .Y(_8418_) );
	OAI21X1 OAI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8418_), .C(_7699_), .Y(_8419_) );
	AOI21X1 AOI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .B(_8041_), .C(_8417_), .Y(_8420_) );
	OAI21X1 OAI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_8043_), .B(_8420_), .C(_8416_), .Y(_8421_) );
	NAND3X1 NAND3X1_1824 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf6), .B(_8421_), .C(_8415_), .Y(_8422_) );
	NAND3X1 NAND3X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf2), .B(_8409_), .C(_8422_), .Y(_8424_) );
	OAI21X1 OAI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_8043_), .B(_8420_), .C(_8410_), .Y(_8425_) );
	NAND3X1 NAND3X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_8416_), .B(_7778_), .C(_8414_), .Y(_8426_) );
	NAND3X1 NAND3X1_1827 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf5), .B(_8425_), .C(_8426_), .Y(_8427_) );
	INVX1 INVX1_1231 ( .gnd(gnd), .vdd(vdd), .A(_8408_), .Y(_8428_) );
	NAND2X1 NAND2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8428_), .B(_8052__bF_buf3), .Y(_8429_) );
	NAND3X1 NAND3X1_1828 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf0), .B(_8429_), .C(_8427_), .Y(_8430_) );
	NAND3X1 NAND3X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .B(_8041_), .C(_8419_), .Y(_8431_) );
	INVX1 INVX1_1232 ( .gnd(gnd), .vdd(vdd), .A(_8431_), .Y(_8432_) );
	OAI21X1 OAI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_8420_), .B(_8432_), .C(divider_divuResult_4_bF_buf4), .Y(_8433_) );
	OAI21X1 OAI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_7668_), .B(_7670_), .C(_8052__bF_buf2), .Y(_8435_) );
	NAND3X1 NAND3X1_1830 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf2), .B(_8435_), .C(_8433_), .Y(_8436_) );
	NAND3X1 NAND3X1_1831 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf3), .B(_8431_), .C(_8414_), .Y(_8437_) );
	INVX1 INVX1_1233 ( .gnd(gnd), .vdd(vdd), .A(_7777_), .Y(_8438_) );
	NAND2X1 NAND2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_8438_), .B(_8052__bF_buf1), .Y(_8439_) );
	NAND3X1 NAND3X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf0), .B(_8439_), .C(_8437_), .Y(_8440_) );
	NAND2X1 NAND2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_8440_), .B(_8436_), .Y(_8441_) );
	NAND3X1 NAND3X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_8424_), .B(_8430_), .C(_8441_), .Y(_8442_) );
	NAND2X1 NAND2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_8037_), .B(_8052__bF_buf0), .Y(_8443_) );
	NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_7765_), .B(_7771_), .Y(_8444_) );
	INVX1 INVX1_1234 ( .gnd(gnd), .vdd(vdd), .A(_8444_), .Y(_8446_) );
	NAND2X1 NAND2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_7697_), .B(_7695_), .Y(_8447_) );
	OAI21X1 OAI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_8418_), .C(_8447_), .Y(_8448_) );
	AOI21X1 AOI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_8448_), .B(_7772_), .C(_8446_), .Y(_8449_) );
	INVX1 INVX1_1235 ( .gnd(gnd), .vdd(vdd), .A(_7693_), .Y(_8450_) );
	OAI21X1 OAI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf0), .B(_8450_), .C(_8448_), .Y(_8451_) );
	NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_8444_), .B(_8451_), .Y(_8452_) );
	OAI21X1 OAI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_8449_), .B(_8452_), .C(divider_divuResult_4_bF_buf2), .Y(_8453_) );
	NAND3X1 NAND3X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf3), .B(_8443_), .C(_8453_), .Y(_8454_) );
	INVX1 INVX1_1236 ( .gnd(gnd), .vdd(vdd), .A(_8037_), .Y(_8455_) );
	NAND2X1 NAND2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_8455_), .B(_8052__bF_buf6), .Y(_8457_) );
	NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_8446_), .B(_8451_), .Y(_8458_) );
	AOI21X1 AOI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_8448_), .B(_7772_), .C(_8444_), .Y(_8459_) );
	OAI21X1 OAI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_8459_), .B(_8458_), .C(divider_divuResult_4_bF_buf1), .Y(_8460_) );
	NAND3X1 NAND3X1_1835 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf3), .B(_8457_), .C(_8460_), .Y(_8461_) );
	INVX1 INVX1_1237 ( .gnd(gnd), .vdd(vdd), .A(_8447_), .Y(_8462_) );
	NAND3X1 NAND3X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_8462_), .B(_7763_), .C(_8411_), .Y(_8463_) );
	NAND2X1 NAND2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_8448_), .B(_8463_), .Y(_8464_) );
	NAND2X1 NAND2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_8464_), .B(divider_divuResult_4_bF_buf0), .Y(_8465_) );
	NAND2X1 NAND2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_8450_), .B(_8052__bF_buf5), .Y(_8466_) );
	NAND3X1 NAND3X1_1837 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .B(_8466_), .C(_8465_), .Y(_8468_) );
	AOI21X1 AOI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_8448_), .B(_8463_), .C(_8052__bF_buf4), .Y(_8469_) );
	INVX1 INVX1_1238 ( .gnd(gnd), .vdd(vdd), .A(_8466_), .Y(_8470_) );
	OAI21X1 OAI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_8470_), .C(_2887__bF_buf1), .Y(_8471_) );
	NAND2X1 NAND2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_8468_), .B(_8471_), .Y(_8472_) );
	NAND3X1 NAND3X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_8454_), .B(_8461_), .C(_8472_), .Y(_8473_) );
	NAND2X1 NAND2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_7759_), .B(_8052__bF_buf3), .Y(_8474_) );
	NAND2X1 NAND2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .B(_7989_), .Y(_8475_) );
	NAND2X1 NAND2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_7994_), .B(_7992_), .Y(_8476_) );
	NAND2X1 NAND2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .B(_8475_), .Y(_8477_) );
	AOI21X1 AOI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7982_), .C(_8477_), .Y(_8479_) );
	OAI21X1 OAI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_7758_), .B(_8479_), .C(_7985_), .Y(_8480_) );
	NAND3X1 NAND3X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_7983_), .B(_7728_), .C(_8480_), .Y(_8481_) );
	OAI21X1 OAI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_8292_), .B(_8289_), .C(_7996_), .Y(_8482_) );
	AOI21X1 AOI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_8482_), .B(_8033_), .C(_7735_), .Y(_8483_) );
	OAI21X1 OAI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_8034_), .B(_8483_), .C(_7724_), .Y(_8484_) );
	NAND3X1 NAND3X1_1840 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf6), .B(_8481_), .C(_8484_), .Y(_8485_) );
	NAND3X1 NAND3X1_1841 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .B(_8474_), .C(_8485_), .Y(_8486_) );
	INVX1 INVX1_1239 ( .gnd(gnd), .vdd(vdd), .A(_7759_), .Y(_8487_) );
	NAND2X1 NAND2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_8487_), .B(_8052__bF_buf2), .Y(_8488_) );
	OAI21X1 OAI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_8034_), .B(_8483_), .C(_7983_), .Y(_8490_) );
	NAND3X1 NAND3X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_7724_), .B(_7728_), .C(_8480_), .Y(_8491_) );
	NAND3X1 NAND3X1_1843 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf5), .B(_8491_), .C(_8490_), .Y(_8492_) );
	NAND3X1 NAND3X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf1), .B(_8488_), .C(_8492_), .Y(_8493_) );
	NAND3X1 NAND3X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_7735_), .B(_8033_), .C(_8482_), .Y(_8494_) );
	NAND2X1 NAND2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_8480_), .B(_8494_), .Y(_8495_) );
	NAND2X1 NAND2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_8495_), .B(divider_divuResult_4_bF_buf4), .Y(_8496_) );
	OAI21X1 OAI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_7732_), .B(divider_divuResult_5_bF_buf3), .C(_7726_), .Y(_8497_) );
	NAND2X1 NAND2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_8497_), .B(_8052__bF_buf1), .Y(_8498_) );
	NAND3X1 NAND3X1_1846 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .B(_8498_), .C(_8496_), .Y(_8499_) );
	AOI21X1 AOI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_8494_), .B(_8480_), .C(_8052__bF_buf0), .Y(_8501_) );
	AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_8052__bF_buf6), .B(_8497_), .Y(_8502_) );
	OAI21X1 OAI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_8501_), .B(_8502_), .C(_1944__bF_buf2), .Y(_8503_) );
	AOI22X1 AOI22X1_184 ( .gnd(gnd), .vdd(vdd), .A(_8499_), .B(_8503_), .C(_8486_), .D(_8493_), .Y(_8504_) );
	INVX1 INVX1_1240 ( .gnd(gnd), .vdd(vdd), .A(_7756_), .Y(_8505_) );
	INVX1 INVX1_1241 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .Y(_8506_) );
	AOI21X1 AOI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_7963_), .B(_7982_), .C(_8506_), .Y(_8507_) );
	OAI21X1 OAI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_8505_), .B(_8507_), .C(_8475_), .Y(_8508_) );
	NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_8505_), .B(_8507_), .Y(_8509_) );
	NAND3X1 NAND3X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .B(_7989_), .C(_8509_), .Y(_8510_) );
	NAND2X1 NAND2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_8508_), .B(_8510_), .Y(_8512_) );
	NAND2X1 NAND2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf3), .B(_8512_), .Y(_8513_) );
	OAI21X1 OAI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_7987_), .B(_7988_), .C(_8052__bF_buf5), .Y(_8514_) );
	NAND3X1 NAND3X1_1848 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf2), .B(_8514_), .C(_8513_), .Y(_8515_) );
	AOI21X1 AOI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_8510_), .B(_8508_), .C(_8052__bF_buf4), .Y(_8516_) );
	AOI21X1 AOI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .B(_7747_), .C(divider_divuResult_4_bF_buf2), .Y(_8517_) );
	OAI21X1 OAI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_8516_), .B(_8517_), .C(_1505__bF_buf0), .Y(_8518_) );
	XNOR2X1 XNOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_8059_), .B(_8506_), .Y(_8519_) );
	OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_8052__bF_buf3), .B(_8519_), .Y(_8520_) );
	NAND3X1 NAND3X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_7754_), .B(_7993_), .C(_8052__bF_buf2), .Y(_8521_) );
	NAND3X1 NAND3X1_1850 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .B(_8521_), .C(_8520_), .Y(_8523_) );
	NAND2X1 NAND2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_8519_), .B(divider_divuResult_4_bF_buf1), .Y(_8524_) );
	NAND2X1 NAND2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_7755_), .B(_8052__bF_buf1), .Y(_8525_) );
	NAND3X1 NAND3X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf2), .B(_8525_), .C(_8524_), .Y(_8526_) );
	AOI22X1 AOI22X1_185 ( .gnd(gnd), .vdd(vdd), .A(_8523_), .B(_8526_), .C(_8518_), .D(_8515_), .Y(_8527_) );
	NAND2X1 NAND2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_8527_), .B(_8504_), .Y(_8528_) );
	NOR3X1 NOR3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_8473_), .B(_8528_), .C(_8442_), .Y(_8529_) );
	NAND3X1 NAND3X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_8407_), .B(_8342_), .C(_8529_), .Y(_8530_) );
	NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_8282_), .B(_8530_), .Y(_8531_) );
	NAND2X1 NAND2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_8407_), .B(_8342_), .Y(_8532_) );
	NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_8473_), .B(_8442_), .Y(_8534_) );
	NAND3X1 NAND3X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf0), .B(_8474_), .C(_8485_), .Y(_8535_) );
	NAND3X1 NAND3X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf4), .B(_8514_), .C(_8513_), .Y(_8536_) );
	AOI21X1 AOI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_8513_), .B(_8514_), .C(_1505__bF_buf3), .Y(_8537_) );
	NAND2X1 NAND2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_8525_), .B(_8524_), .Y(_8538_) );
	NAND2X1 NAND2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf1), .B(_8538_), .Y(_8539_) );
	AOI21X1 AOI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .B(_8536_), .C(_8537_), .Y(_8540_) );
	NAND2X1 NAND2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_8504_), .B(_8540_), .Y(_8541_) );
	OAI21X1 OAI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_8487_), .B(divider_divuResult_4_bF_buf0), .C(_8485_), .Y(_8542_) );
	INVX1 INVX1_1242 ( .gnd(gnd), .vdd(vdd), .A(_8542_), .Y(_8543_) );
	NAND3X1 NAND3X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf1), .B(_8498_), .C(_8496_), .Y(_8545_) );
	INVX1 INVX1_1243 ( .gnd(gnd), .vdd(vdd), .A(_8545_), .Y(_8546_) );
	OAI21X1 OAI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf3), .B(_8543_), .C(_8546_), .Y(_8547_) );
	NAND3X1 NAND3X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_8535_), .B(_8547_), .C(_8541_), .Y(_8548_) );
	AOI21X1 AOI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_8460_), .B(_8457_), .C(divider_absoluteValue_B_flipSign_result_18_bF_buf2), .Y(_8549_) );
	OAI21X1 OAI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_7693_), .B(divider_divuResult_4_bF_buf6), .C(_8465_), .Y(_8550_) );
	NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .B(_8550_), .Y(_8551_) );
	AOI21X1 AOI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_8551_), .B(_8461_), .C(_8549_), .Y(_8552_) );
	AOI21X1 AOI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_8427_), .B(_8429_), .C(divider_absoluteValue_B_flipSign_result_20_bF_buf3), .Y(_8553_) );
	NAND3X1 NAND3X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf4), .B(_8435_), .C(_8433_), .Y(_8554_) );
	INVX1 INVX1_1244 ( .gnd(gnd), .vdd(vdd), .A(_8554_), .Y(_8556_) );
	AOI21X1 AOI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_8556_), .B(_8430_), .C(_8553_), .Y(_8557_) );
	OAI21X1 OAI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_8552_), .B(_8442_), .C(_8557_), .Y(_8558_) );
	AOI21X1 AOI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_8548_), .B(_8534_), .C(_8558_), .Y(_8559_) );
	OAI21X1 OAI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_8399_), .B(_8403_), .C(divider_absoluteValue_B_flipSign_result_22_bF_buf3), .Y(_8560_) );
	OAI21X1 OAI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_7597_), .B(divider_divuResult_4_bF_buf5), .C(_8383_), .Y(_8561_) );
	NAND3X1 NAND3X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf0), .B(_8392_), .C(_8397_), .Y(_8562_) );
	OAI21X1 OAI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf0), .B(_8561_), .C(_8562_), .Y(_8563_) );
	NAND2X1 NAND2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_8560_), .B(_8563_), .Y(_8564_) );
	AOI21X1 AOI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_8362_), .B(_8364_), .C(divider_absoluteValue_B_flipSign_result_24_bF_buf0), .Y(_8565_) );
	NAND3X1 NAND3X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf0), .B(_8370_), .C(_8369_), .Y(_8567_) );
	INVX1 INVX1_1245 ( .gnd(gnd), .vdd(vdd), .A(_8567_), .Y(_8568_) );
	AOI21X1 AOI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_8568_), .B(_8365_), .C(_8565_), .Y(_8569_) );
	OAI21X1 OAI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_8564_), .B(_8377_), .C(_8569_), .Y(_8570_) );
	NOR3X1 NOR3X1_85 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf1), .B(_8326_), .C(_8329_), .Y(_8571_) );
	NAND2X1 NAND2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_8338_), .B(_8337_), .Y(_8572_) );
	NAND2X1 NAND2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_8572_), .Y(_8573_) );
	INVX1 INVX1_1246 ( .gnd(gnd), .vdd(vdd), .A(_8573_), .Y(_8574_) );
	AOI21X1 AOI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_8330_), .B(_8574_), .C(_8571_), .Y(_8575_) );
	NAND2X1 NAND2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_8283_), .Y(_8576_) );
	INVX1 INVX1_1247 ( .gnd(gnd), .vdd(vdd), .A(_8576_), .Y(_8578_) );
	AOI21X1 AOI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_8311_), .B(_8312_), .C(divider_absoluteValue_B_flipSign_result_27_), .Y(_8579_) );
	AOI21X1 AOI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_8579_), .B(_8286_), .C(_8578_), .Y(_8580_) );
	OAI21X1 OAI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8575_), .C(_8580_), .Y(_8581_) );
	AOI21X1 AOI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_8342_), .B(_8570_), .C(_8581_), .Y(_8582_) );
	OAI21X1 OAI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_8532_), .B(_8559_), .C(_8582_), .Y(_8583_) );
	NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf4), .B(_1571_), .Y(_8584_) );
	OAI21X1 OAI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_8531_), .B(_8583_), .C(_8584_), .Y(_8585_) );
	NAND2X1 NAND2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_3_), .B(_8585_), .Y(_8586_) );
	INVX1 INVX1_1248 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_3_), .Y(_8587_) );
	NAND3X1 NAND3X1_1860 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf3), .B(_8344_), .C(_8358_), .Y(_8589_) );
	NAND3X1 NAND3X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf2), .B(_8364_), .C(_8362_), .Y(_8590_) );
	NAND2X1 NAND2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_8589_), .B(_8590_), .Y(_8591_) );
	AOI22X1 AOI22X1_186 ( .gnd(gnd), .vdd(vdd), .A(_8385_), .B(_8389_), .C(_8398_), .D(_8404_), .Y(_8592_) );
	NAND3X1 NAND3X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_8376_), .B(_8592_), .C(_8591_), .Y(_8593_) );
	NOR3X1 NOR3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_8341_), .C(_8593_), .Y(_8594_) );
	AOI21X1 AOI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_8018_), .B(_8053_), .C(_1735__bF_buf6), .Y(_8595_) );
	OAI21X1 OAI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_8074_), .B(divider_divuResult_4_bF_buf4), .C(_8077_), .Y(_8596_) );
	NAND2X1 NAND2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_8596_), .Y(_8597_) );
	OAI21X1 OAI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_8597_), .B(_8595_), .C(_8054_), .Y(_8598_) );
	NAND3X1 NAND3X1_1863 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_8105_), .C(_8103_), .Y(_8600_) );
	NAND3X1 NAND3X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_8090_), .C(_8600_), .Y(_8601_) );
	NAND2X1 NAND2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_8105_), .B(_8103_), .Y(_8602_) );
	AOI22X1 AOI22X1_187 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_2547__bF_buf0), .C(_1768__bF_buf7), .D(_8602_), .Y(_8603_) );
	AOI21X1 AOI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_8601_), .B(_8603_), .C(_8087_), .Y(_8604_) );
	AOI21X1 AOI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_8604_), .B(_8080_), .C(_8598_), .Y(_8605_) );
	AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_8171_), .B(_8200_), .Y(_8606_) );
	AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_8271_), .B(_8253_), .Y(_8607_) );
	NAND2X1 NAND2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_8607_), .B(_8606_), .Y(_8608_) );
	OAI21X1 OAI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_8151_), .B(_8150_), .C(_1484__bF_buf3), .Y(_8609_) );
	NAND2X1 NAND2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_8164_), .B(_8169_), .Y(_8611_) );
	NAND3X1 NAND3X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_8256_), .B(_8609_), .C(_8611_), .Y(_8612_) );
	INVX1 INVX1_1249 ( .gnd(gnd), .vdd(vdd), .A(_8609_), .Y(_8613_) );
	AOI21X1 AOI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_8166_), .B(_8168_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf2), .Y(_8614_) );
	OAI21X1 OAI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(_8613_), .C(_8256_), .Y(_8615_) );
	OAI21X1 OAI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_8182_), .B(divider_divuResult_4_bF_buf3), .C(_8179_), .Y(_8616_) );
	INVX1 INVX1_1250 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .Y(_8617_) );
	OAI21X1 OAI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_8197_), .B(divider_divuResult_4_bF_buf2), .C(_8193_), .Y(_8618_) );
	OAI21X1 OAI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf1), .B(_8618_), .C(_8265_), .Y(_8619_) );
	OAI21X1 OAI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf4), .B(_8617_), .C(_8619_), .Y(_8620_) );
	OAI21X1 OAI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_8620_), .B(_8612_), .C(_8615_), .Y(_8622_) );
	NOR3X1 NOR3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf4), .B(_8212_), .C(_8213_), .Y(_8623_) );
	AOI21X1 AOI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_8210_), .B(_8202_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .Y(_8624_) );
	OAI21X1 OAI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_8624_), .B(_8623_), .C(_8228_), .Y(_8625_) );
	NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_8212_), .B(_8213_), .Y(_8626_) );
	OAI21X1 OAI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf3), .B(_8626_), .C(_8274_), .Y(_8627_) );
	OAI21X1 OAI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_8239_), .B(divider_divuResult_4_bF_buf1), .C(_8237_), .Y(_8628_) );
	NAND2X1 NAND2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_8628_), .Y(_8629_) );
	OAI21X1 OAI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .B(divider_divuResult_4_bF_buf0), .C(_8246_), .Y(_8630_) );
	OAI21X1 OAI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf6), .B(_8630_), .C(_8275_), .Y(_8631_) );
	NAND2X1 NAND2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_8629_), .B(_8631_), .Y(_8633_) );
	OAI21X1 OAI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_8633_), .B(_8625_), .C(_8627_), .Y(_8634_) );
	AOI21X1 AOI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_8634_), .B(_8606_), .C(_8622_), .Y(_8635_) );
	OAI21X1 OAI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_8605_), .B(_8608_), .C(_8635_), .Y(_8636_) );
	NAND3X1 NAND3X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_8529_), .B(_8594_), .C(_8636_), .Y(_8637_) );
	NAND3X1 NAND3X1_1867 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf2), .B(_8409_), .C(_8422_), .Y(_8638_) );
	NAND3X1 NAND3X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf1), .B(_8429_), .C(_8427_), .Y(_8639_) );
	AOI22X1 AOI22X1_188 ( .gnd(gnd), .vdd(vdd), .A(_8436_), .B(_8440_), .C(_8638_), .D(_8639_), .Y(_8640_) );
	NAND3X1 NAND3X1_1869 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf1), .B(_8443_), .C(_8453_), .Y(_8641_) );
	NAND3X1 NAND3X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf2), .B(_8457_), .C(_8460_), .Y(_8642_) );
	AOI22X1 AOI22X1_189 ( .gnd(gnd), .vdd(vdd), .A(_8468_), .B(_8471_), .C(_8642_), .D(_8641_), .Y(_8644_) );
	NAND2X1 NAND2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .B(_8640_), .Y(_8645_) );
	AOI21X1 AOI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_8485_), .B(_8474_), .C(_2922__bF_buf2), .Y(_8646_) );
	OAI21X1 OAI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_8545_), .B(_8646_), .C(_8535_), .Y(_8647_) );
	AOI21X1 AOI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_8540_), .B(_8504_), .C(_8647_), .Y(_8648_) );
	AOI21X1 AOI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_8453_), .B(_8443_), .C(_3263__bF_buf1), .Y(_8649_) );
	NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_8470_), .Y(_8650_) );
	NAND2X1 NAND2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf0), .B(_8650_), .Y(_8651_) );
	OAI21X1 OAI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8649_), .C(_8454_), .Y(_8652_) );
	AOI21X1 AOI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_8422_), .B(_8409_), .C(_4011__bF_buf0), .Y(_8653_) );
	OAI21X1 OAI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_8554_), .B(_8653_), .C(_8424_), .Y(_8655_) );
	AOI21X1 AOI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8652_), .C(_8655_), .Y(_8656_) );
	OAI21X1 OAI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_8645_), .B(_8648_), .C(_8656_), .Y(_8657_) );
	NAND2X1 NAND2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_8594_), .B(_8657_), .Y(_8658_) );
	NAND3X1 NAND3X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_8582_), .B(_8658_), .C(_8637_), .Y(_8659_) );
	NAND3X1 NAND3X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_8587_), .B(_8584_), .C(_8659_), .Y(_8660_) );
	NAND2X1 NAND2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_8660_), .B(_8586_), .Y(_8661_) );
	NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_30_), .B(divider_absoluteValue_B_flipSign_result_31_), .Y(_8662_) );
	INVX1 INVX1_1251 ( .gnd(gnd), .vdd(vdd), .A(_8662_), .Y(_8663_) );
	OAI21X1 OAI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_8531_), .B(_8583_), .C(_2020_), .Y(_8664_) );
	AOI21X1 AOI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_8664__bF_buf6), .B(_8283_), .C(_2240__bF_buf4), .Y(_8666_) );
	INVX1 INVX1_1252 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .Y(_8667_) );
	NAND2X1 NAND2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .B(_8667_), .Y(_8668_) );
	NAND2X1 NAND2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_8666_), .Y(_8669_) );
	NAND3X1 NAND3X1_1873 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_8306_), .C(_8304_), .Y(_8670_) );
	NAND3X1 NAND3X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_8312_), .C(_8311_), .Y(_8671_) );
	AOI22X1 AOI22X1_190 ( .gnd(gnd), .vdd(vdd), .A(_8284_), .B(_8285_), .C(_8671_), .D(_8670_), .Y(_8672_) );
	NAND3X1 NAND3X1_1875 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf0), .B(_8316_), .C(_8323_), .Y(_8673_) );
	OAI21X1 OAI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_8326_), .B(_8329_), .C(_6845_), .Y(_8674_) );
	AOI22X1 AOI22X1_191 ( .gnd(gnd), .vdd(vdd), .A(_8336_), .B(_8339_), .C(_8673_), .D(_8674_), .Y(_8675_) );
	NAND2X1 NAND2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_8672_), .B(_8675_), .Y(_8677_) );
	AOI22X1 AOI22X1_192 ( .gnd(gnd), .vdd(vdd), .A(_8371_), .B(_8375_), .C(_8589_), .D(_8590_), .Y(_8678_) );
	AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_8563_), .B(_8560_), .Y(_8679_) );
	AOI21X1 AOI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_8358_), .B(_8344_), .C(_2042__bF_buf1), .Y(_8680_) );
	OAI21X1 OAI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_8567_), .B(_8680_), .C(_8359_), .Y(_8681_) );
	AOI21X1 AOI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_8679_), .B(_8678_), .C(_8681_), .Y(_8682_) );
	AOI21X1 AOI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_8323_), .B(_8316_), .C(_6845_), .Y(_8683_) );
	OAI21X1 OAI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_8573_), .B(_8683_), .C(_8325_), .Y(_8684_) );
	NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_8283_), .Y(_8685_) );
	OAI21X1 OAI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_8685_), .B(_8307_), .C(_8576_), .Y(_8686_) );
	AOI21X1 AOI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_8672_), .B(_8684_), .C(_8686_), .Y(_8688_) );
	OAI21X1 OAI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_8677_), .B(_8682_), .C(_8688_), .Y(_8689_) );
	AOI21X1 AOI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_8594_), .B(_8657_), .C(_8689_), .Y(_8690_) );
	AOI21X1 AOI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_8690_), .B(_8637_), .C(_1571_), .Y(divider_divuResult_3_) );
	AOI21X1 AOI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_8080_), .B(_8095_), .C(_8598_), .Y(_8691_) );
	AOI21X1 AOI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_8691_), .B(_8112_), .C(_8608_), .Y(_8692_) );
	OAI21X1 OAI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .B(_8692_), .C(_8529_), .Y(_8693_) );
	AOI21X1 AOI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_8693_), .B(_8559_), .C(_8593_), .Y(_8694_) );
	OAI21X1 OAI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_8570_), .B(_8694_), .C(_8675_), .Y(_8695_) );
	AOI22X1 AOI22X1_193 ( .gnd(gnd), .vdd(vdd), .A(_8670_), .B(_8671_), .C(_8575_), .D(_8695_), .Y(_8696_) );
	NAND2X1 NAND2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_8671_), .B(_8670_), .Y(_8698_) );
	NAND2X1 NAND2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_8255_), .B(_8113_), .Y(_8699_) );
	INVX1 INVX1_1253 ( .gnd(gnd), .vdd(vdd), .A(_8528_), .Y(_8700_) );
	NAND3X1 NAND3X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .B(_8640_), .C(_8700_), .Y(_8701_) );
	AOI21X1 AOI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_8699_), .B(_8635_), .C(_8701_), .Y(_8702_) );
	OAI21X1 OAI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_8657_), .B(_8702_), .C(_8407_), .Y(_8703_) );
	AOI21X1 AOI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_8703_), .B(_8682_), .C(_8341_), .Y(_8704_) );
	NOR3X1 NOR3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_8698_), .B(_8684_), .C(_8704_), .Y(_8705_) );
	OAI21X1 OAI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_8696_), .B(_8705_), .C(divider_divuResult_3_bF_buf7), .Y(_8706_) );
	OAI21X1 OAI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_8305_), .B(divider_divuResult_4_bF_buf6), .C(_8304_), .Y(_8707_) );
	NAND2X1 NAND2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_8707_), .B(_8664__bF_buf5), .Y(_8709_) );
	NAND3X1 NAND3X1_1877 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .B(_8709_), .C(_8706_), .Y(_8710_) );
	OAI21X1 OAI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .B(_8704_), .C(_8698_), .Y(_8711_) );
	INVX1 INVX1_1254 ( .gnd(gnd), .vdd(vdd), .A(_8698_), .Y(_8712_) );
	NAND3X1 NAND3X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_8712_), .B(_8575_), .C(_8695_), .Y(_8713_) );
	NAND3X1 NAND3X1_1879 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf6), .B(_8711_), .C(_8713_), .Y(_8714_) );
	OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf5), .B(_8707_), .Y(_8715_) );
	NAND3X1 NAND3X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_8715_), .C(_8714_), .Y(_8716_) );
	AOI22X1 AOI22X1_194 ( .gnd(gnd), .vdd(vdd), .A(_8668_), .B(_8669_), .C(_8716_), .D(_8710_), .Y(_8717_) );
	OAI21X1 OAI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_8326_), .B(_8329_), .C(_8664__bF_buf4), .Y(_8718_) );
	NAND2X1 NAND2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_8673_), .B(_8674_), .Y(_8720_) );
	OAI21X1 OAI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_8570_), .B(_8694_), .C(_8340_), .Y(_8721_) );
	NAND3X1 NAND3X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_8720_), .B(_8573_), .C(_8721_), .Y(_8722_) );
	INVX1 INVX1_1255 ( .gnd(gnd), .vdd(vdd), .A(_8720_), .Y(_8723_) );
	INVX1 INVX1_1256 ( .gnd(gnd), .vdd(vdd), .A(_8340_), .Y(_8724_) );
	AOI21X1 AOI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_8703_), .B(_8682_), .C(_8724_), .Y(_8725_) );
	OAI21X1 OAI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_8574_), .B(_8725_), .C(_8723_), .Y(_8726_) );
	NAND3X1 NAND3X1_1882 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf4), .B(_8726_), .C(_8722_), .Y(_8727_) );
	NAND3X1 NAND3X1_1883 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_8718_), .C(_8727_), .Y(_8728_) );
	INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(_8718_), .Y(_8729_) );
	OAI21X1 OAI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_8574_), .B(_8725_), .C(_8720_), .Y(_8730_) );
	NAND3X1 NAND3X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_8723_), .B(_8573_), .C(_8721_), .Y(_8731_) );
	AOI21X1 AOI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_8731_), .B(_8730_), .C(_8664__bF_buf3), .Y(_8732_) );
	OAI21X1 OAI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_8729_), .B(_8732_), .C(_7453_), .Y(_8733_) );
	OAI21X1 OAI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_8701_), .B(_8282_), .C(_8559_), .Y(_8734_) );
	AOI21X1 AOI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .B(_8407_), .C(_8570_), .Y(_8735_) );
	AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8724_), .Y(_8736_) );
	OAI21X1 OAI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_8724_), .B(_8735_), .C(divider_divuResult_3_bF_buf3), .Y(_8737_) );
	NAND2X1 NAND2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_8572_), .B(_8664__bF_buf2), .Y(_8738_) );
	OAI21X1 OAI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_8737_), .C(_8738_), .Y(_8739_) );
	XNOR2X1 XNOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_6845_), .Y(_8741_) );
	AOI21X1 AOI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_8733_), .B(_8728_), .C(_8741_), .Y(_8742_) );
	NAND2X1 NAND2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_8717_), .B(_8742_), .Y(_8743_) );
	OAI21X1 OAI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_8363_), .B(divider_divuResult_4_bF_buf5), .C(_8358_), .Y(_8744_) );
	NAND2X1 NAND2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_8744_), .B(_8664__bF_buf1), .Y(_8745_) );
	AOI21X1 AOI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_8693_), .B(_8559_), .C(_8406_), .Y(_8746_) );
	OAI21X1 OAI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_8679_), .B(_8746_), .C(_8376_), .Y(_8747_) );
	NAND3X1 NAND3X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_8567_), .C(_8747_), .Y(_8748_) );
	INVX1 INVX1_1257 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .Y(_8749_) );
	OAI21X1 OAI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_8657_), .B(_8702_), .C(_8592_), .Y(_8750_) );
	AOI22X1 AOI22X1_195 ( .gnd(gnd), .vdd(vdd), .A(_8371_), .B(_8375_), .C(_8564_), .D(_8750_), .Y(_8752_) );
	OAI21X1 OAI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_8568_), .B(_8752_), .C(_8749_), .Y(_8753_) );
	NAND3X1 NAND3X1_1886 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf2), .B(_8753_), .C(_8748_), .Y(_8754_) );
	NAND3X1 NAND3X1_1887 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_8745_), .C(_8754_), .Y(_8755_) );
	INVX1 INVX1_1258 ( .gnd(gnd), .vdd(vdd), .A(_8744_), .Y(_8756_) );
	NAND2X1 NAND2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_8756_), .B(_8664__bF_buf0), .Y(_8757_) );
	OAI21X1 OAI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_8568_), .B(_8752_), .C(_8591_), .Y(_8758_) );
	NAND3X1 NAND3X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_8749_), .B(_8567_), .C(_8747_), .Y(_8759_) );
	NAND3X1 NAND3X1_1889 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf1), .B(_8758_), .C(_8759_), .Y(_8760_) );
	NAND3X1 NAND3X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_8757_), .C(_8760_), .Y(_8761_) );
	INVX1 INVX1_1259 ( .gnd(gnd), .vdd(vdd), .A(_8376_), .Y(_8763_) );
	NAND3X1 NAND3X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_8763_), .B(_8564_), .C(_8750_), .Y(_8764_) );
	INVX1 INVX1_1260 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .Y(_8765_) );
	OAI21X1 OAI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_8752_), .B(_8765_), .C(divider_divuResult_3_bF_buf0), .Y(_8766_) );
	OAI21X1 OAI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .B(_8374_), .C(_8664__bF_buf6), .Y(_8767_) );
	NAND3X1 NAND3X1_1892 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf2), .B(_8767_), .C(_8766_), .Y(_8768_) );
	AOI21X1 AOI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_8747_), .B(_8764_), .C(_8664__bF_buf5), .Y(_8769_) );
	OAI21X1 OAI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_8373_), .B(divider_divuResult_4_bF_buf4), .C(_8369_), .Y(_8770_) );
	INVX1 INVX1_1261 ( .gnd(gnd), .vdd(vdd), .A(_8770_), .Y(_8771_) );
	NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(divider_divuResult_3_bF_buf7), .Y(_8772_) );
	OAI21X1 OAI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_8772_), .B(_8769_), .C(_2042__bF_buf0), .Y(_8774_) );
	AOI22X1 AOI22X1_196 ( .gnd(gnd), .vdd(vdd), .A(_8768_), .B(_8774_), .C(_8755_), .D(_8761_), .Y(_8775_) );
	OAI21X1 OAI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_8399_), .B(_8403_), .C(_8664__bF_buf4), .Y(_8776_) );
	INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(_8776_), .Y(_8777_) );
	INVX1 INVX1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8561_), .Y(_8778_) );
	NAND2X1 NAND2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf0), .B(_8778_), .Y(_8779_) );
	OAI21X1 OAI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_8657_), .B(_8702_), .C(_8391_), .Y(_8780_) );
	NAND3X1 NAND3X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_8405_), .C(_8780_), .Y(_8781_) );
	INVX1 INVX1_1263 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .Y(_8782_) );
	INVX1 INVX1_1264 ( .gnd(gnd), .vdd(vdd), .A(_8405_), .Y(_8783_) );
	INVX1 INVX1_1265 ( .gnd(gnd), .vdd(vdd), .A(_8391_), .Y(_8785_) );
	AOI21X1 AOI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_8693_), .B(_8559_), .C(_8785_), .Y(_8786_) );
	OAI21X1 OAI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .B(_8786_), .C(_8783_), .Y(_8787_) );
	NAND3X1 NAND3X1_1894 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf6), .B(_8781_), .C(_8787_), .Y(_8788_) );
	INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(_8788_), .Y(_8789_) );
	OAI21X1 OAI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_8777_), .B(_8789_), .C(divider_absoluteValue_B_flipSign_result_23_bF_buf0), .Y(_8790_) );
	NAND3X1 NAND3X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf3), .B(_8776_), .C(_8788_), .Y(_8791_) );
	NAND3X1 NAND3X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8559_), .C(_8693_), .Y(_8792_) );
	INVX1 INVX1_1266 ( .gnd(gnd), .vdd(vdd), .A(_8792_), .Y(_8793_) );
	OAI21X1 OAI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_8786_), .B(_8793_), .C(divider_divuResult_3_bF_buf5), .Y(_8794_) );
	OAI21X1 OAI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_8778_), .B(divider_divuResult_3_bF_buf4), .C(_8794_), .Y(_8796_) );
	OAI21X1 OAI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf2), .B(_8796_), .C(_8791_), .Y(_8797_) );
	AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_8797_), .B(_8790_), .Y(_8798_) );
	NAND3X1 NAND3X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_8745_), .C(_8754_), .Y(_8799_) );
	AOI21X1 AOI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_8754_), .B(_8745_), .C(_2053_), .Y(_8800_) );
	NAND3X1 NAND3X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf3), .B(_8767_), .C(_8766_), .Y(_8801_) );
	OAI21X1 OAI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_8801_), .B(_8800_), .C(_8799_), .Y(_8802_) );
	AOI21X1 AOI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_8775_), .B(_8798_), .C(_8802_), .Y(_8803_) );
	NAND3X1 NAND3X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_8718_), .C(_8727_), .Y(_8804_) );
	AOI21X1 AOI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_8727_), .B(_8718_), .C(_7453_), .Y(_8805_) );
	NAND2X1 NAND2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_8739_), .Y(_8807_) );
	OAI21X1 OAI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_8807_), .B(_8805_), .C(_8804_), .Y(_8808_) );
	NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .B(_8666_), .Y(_8809_) );
	INVX1 INVX1_1267 ( .gnd(gnd), .vdd(vdd), .A(_8809_), .Y(_8810_) );
	NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_8667_), .Y(_8811_) );
	NAND3X1 NAND3X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_8709_), .C(_8706_), .Y(_8812_) );
	OAI21X1 OAI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8812_), .C(_8810_), .Y(_8813_) );
	AOI21X1 AOI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_8717_), .B(_8808_), .C(_8813_), .Y(_8814_) );
	OAI21X1 OAI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_8803_), .B(_8743_), .C(_8814_), .Y(_8815_) );
	NAND2X1 NAND2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_8669_), .B(_8668_), .Y(_8816_) );
	NAND3X1 NAND3X1_1901 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .B(_8715_), .C(_8714_), .Y(_8818_) );
	NAND3X1 NAND3X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8818_), .C(_8812_), .Y(_8819_) );
	OAI21X1 OAI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_8729_), .B(_8732_), .C(divider_absoluteValue_B_flipSign_result_27_), .Y(_8820_) );
	XNOR2X1 XNOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(divider_absoluteValue_B_flipSign_result_26_bF_buf3), .Y(_8821_) );
	NAND3X1 NAND3X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_8804_), .B(_8820_), .C(_8821_), .Y(_8822_) );
	NAND3X1 NAND3X1_1904 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf3), .B(_8776_), .C(_8788_), .Y(_8823_) );
	OAI21X1 OAI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_8777_), .B(_8789_), .C(_5516__bF_buf2), .Y(_8824_) );
	OAI21X1 OAI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_8387_), .B(_8388_), .C(_8664__bF_buf3), .Y(_8825_) );
	NAND3X1 NAND3X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf3), .B(_8825_), .C(_8794_), .Y(_8826_) );
	NAND2X1 NAND2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf1), .B(_8796_), .Y(_8827_) );
	NAND2X1 NAND2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_8826_), .B(_8827_), .Y(_8829_) );
	AOI21X1 AOI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_8824_), .B(_8823_), .C(_8829_), .Y(_8830_) );
	NAND2X1 NAND2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_8830_), .B(_8775_), .Y(_8831_) );
	NOR3X1 NOR3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_8819_), .B(_8822_), .C(_8831_), .Y(_8832_) );
	OAI21X1 OAI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_8428_), .B(divider_divuResult_4_bF_buf3), .C(_8422_), .Y(_8833_) );
	NAND2X1 NAND2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_8833_), .B(_8664__bF_buf2), .Y(_8834_) );
	NAND2X1 NAND2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_8638_), .B(_8639_), .Y(_8835_) );
	OAI21X1 OAI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .B(_8692_), .C(_8700_), .Y(_8836_) );
	AOI21X1 AOI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_8836_), .B(_8648_), .C(_8473_), .Y(_8837_) );
	OAI21X1 OAI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_8652_), .B(_8837_), .C(_8441_), .Y(_8838_) );
	NAND3X1 NAND3X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_8554_), .C(_8838_), .Y(_8840_) );
	INVX1 INVX1_1268 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .Y(_8841_) );
	INVX1 INVX1_1269 ( .gnd(gnd), .vdd(vdd), .A(_8441_), .Y(_8842_) );
	AOI21X1 AOI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_8699_), .B(_8635_), .C(_8528_), .Y(_8843_) );
	OAI21X1 OAI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_8548_), .B(_8843_), .C(_8644_), .Y(_8844_) );
	AOI21X1 AOI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_8844_), .B(_8552_), .C(_8842_), .Y(_8845_) );
	OAI21X1 OAI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_8556_), .B(_8845_), .C(_8841_), .Y(_8846_) );
	NAND3X1 NAND3X1_1907 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf3), .B(_8846_), .C(_8840_), .Y(_8847_) );
	NAND3X1 NAND3X1_1908 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf3), .B(_8834_), .C(_8847_), .Y(_8848_) );
	INVX1 INVX1_1270 ( .gnd(gnd), .vdd(vdd), .A(_8833_), .Y(_8849_) );
	NAND2X1 NAND2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_8849_), .B(_8664__bF_buf1), .Y(_8851_) );
	OAI21X1 OAI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_8556_), .B(_8845_), .C(_8835_), .Y(_8852_) );
	NAND3X1 NAND3X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_8554_), .C(_8838_), .Y(_8853_) );
	NAND3X1 NAND3X1_1910 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf2), .B(_8852_), .C(_8853_), .Y(_8854_) );
	NAND3X1 NAND3X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf3), .B(_8851_), .C(_8854_), .Y(_8855_) );
	OAI21X1 OAI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_8528_), .B(_8282_), .C(_8648_), .Y(_8856_) );
	AOI21X1 AOI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_8856_), .B(_8644_), .C(_8652_), .Y(_8857_) );
	AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_8842_), .Y(_8858_) );
	OAI21X1 OAI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_8858_), .C(divider_divuResult_3_bF_buf1), .Y(_8859_) );
	OAI21X1 OAI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_8438_), .B(divider_divuResult_4_bF_buf2), .C(_8433_), .Y(_8860_) );
	NAND2X1 NAND2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_8664__bF_buf0), .Y(_8862_) );
	NAND3X1 NAND3X1_1912 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf1), .B(_8862_), .C(_8859_), .Y(_8863_) );
	NAND2X1 NAND2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_8842_), .B(_8857_), .Y(_8864_) );
	NAND3X1 NAND3X1_1913 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf0), .B(_8864_), .C(_8838_), .Y(_8865_) );
	OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf7), .B(_8860_), .Y(_8866_) );
	NAND3X1 NAND3X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf3), .B(_8866_), .C(_8865_), .Y(_8867_) );
	AOI22X1 AOI22X1_197 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .B(_8867_), .C(_8848_), .D(_8855_), .Y(_8868_) );
	OAI21X1 OAI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_8455_), .B(divider_divuResult_4_bF_buf1), .C(_8453_), .Y(_8869_) );
	NAND2X1 NAND2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_8869_), .B(_8664__bF_buf6), .Y(_8870_) );
	NAND2X1 NAND2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_8642_), .B(_8641_), .Y(_8871_) );
	OAI21X1 OAI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_8548_), .B(_8843_), .C(_8472_), .Y(_8873_) );
	OAI21X1 OAI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .B(_8550_), .C(_8873_), .Y(_8874_) );
	AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_8874_), .B(_8871_), .Y(_8875_) );
	NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8874_), .Y(_8876_) );
	OAI21X1 OAI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_8876_), .B(_8875_), .C(divider_divuResult_3_bF_buf6), .Y(_8877_) );
	NAND3X1 NAND3X1_1915 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf1), .B(_8870_), .C(_8877_), .Y(_8878_) );
	INVX1 INVX1_1271 ( .gnd(gnd), .vdd(vdd), .A(_8869_), .Y(_8879_) );
	NAND2X1 NAND2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_8664__bF_buf5), .Y(_8880_) );
	NAND2X1 NAND2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8874_), .Y(_8881_) );
	OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_8874_), .B(_8871_), .Y(_8882_) );
	NAND3X1 NAND3X1_1916 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf5), .B(_8881_), .C(_8882_), .Y(_8884_) );
	NAND3X1 NAND3X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf3), .B(_8880_), .C(_8884_), .Y(_8885_) );
	OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_8856_), .B(_8472_), .Y(_8886_) );
	NAND2X1 NAND2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_8873_), .B(_8886_), .Y(_8887_) );
	NAND2X1 NAND2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf4), .B(_8887_), .Y(_8888_) );
	OAI21X1 OAI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_8470_), .C(_8664__bF_buf4), .Y(_8889_) );
	NAND3X1 NAND3X1_1918 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf0), .B(_8889_), .C(_8888_), .Y(_8890_) );
	NAND3X1 NAND3X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_8873_), .B(_8886_), .C(divider_divuResult_3_bF_buf3), .Y(_8891_) );
	NAND2X1 NAND2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_8650_), .B(_8664__bF_buf3), .Y(_8892_) );
	NAND3X1 NAND3X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf0), .B(_8892_), .C(_8891_), .Y(_8893_) );
	AOI22X1 AOI22X1_198 ( .gnd(gnd), .vdd(vdd), .A(_8890_), .B(_8893_), .C(_8885_), .D(_8878_), .Y(_8895_) );
	NAND2X1 NAND2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_8895_), .B(_8868_), .Y(_8896_) );
	NAND2X1 NAND2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_8542_), .B(_8664__bF_buf2), .Y(_8897_) );
	NAND2X1 NAND2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .B(_8493_), .Y(_8898_) );
	NAND2X1 NAND2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_8499_), .B(_8503_), .Y(_8899_) );
	INVX1 INVX1_1272 ( .gnd(gnd), .vdd(vdd), .A(_8527_), .Y(_8900_) );
	INVX1 INVX1_1273 ( .gnd(gnd), .vdd(vdd), .A(_8540_), .Y(_8901_) );
	OAI21X1 OAI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_8900_), .B(_8282_), .C(_8901_), .Y(_8902_) );
	NAND2X1 NAND2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_8899_), .B(_8902_), .Y(_8903_) );
	NAND3X1 NAND3X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_8898_), .B(_8545_), .C(_8903_), .Y(_8904_) );
	INVX1 INVX1_1274 ( .gnd(gnd), .vdd(vdd), .A(_8898_), .Y(_8906_) );
	INVX1 INVX1_1275 ( .gnd(gnd), .vdd(vdd), .A(_8899_), .Y(_8907_) );
	OAI21X1 OAI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .B(_8692_), .C(_8527_), .Y(_8908_) );
	AOI21X1 AOI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8901_), .C(_8907_), .Y(_8909_) );
	OAI21X1 OAI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_8546_), .B(_8909_), .C(_8906_), .Y(_8910_) );
	NAND3X1 NAND3X1_1922 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf2), .B(_8904_), .C(_8910_), .Y(_8911_) );
	NAND3X1 NAND3X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf4), .B(_8897_), .C(_8911_), .Y(_8912_) );
	NAND2X1 NAND2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_8543_), .B(_8664__bF_buf1), .Y(_8913_) );
	OAI21X1 OAI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_8546_), .B(_8909_), .C(_8898_), .Y(_8914_) );
	NAND3X1 NAND3X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_8906_), .B(_8545_), .C(_8903_), .Y(_8915_) );
	NAND3X1 NAND3X1_1925 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf1), .B(_8915_), .C(_8914_), .Y(_8917_) );
	NAND3X1 NAND3X1_1926 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf0), .B(_8913_), .C(_8917_), .Y(_8918_) );
	NAND2X1 NAND2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_8912_), .B(_8918_), .Y(_8919_) );
	NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_8899_), .B(_8902_), .Y(_8920_) );
	OAI21X1 OAI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_8920_), .C(divider_divuResult_3_bF_buf0), .Y(_8921_) );
	OAI21X1 OAI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_8501_), .B(_8502_), .C(_8664__bF_buf0), .Y(_8922_) );
	NAND3X1 NAND3X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_2922__bF_buf1), .B(_8921_), .C(_8922_), .Y(_8923_) );
	NAND3X1 NAND3X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8901_), .C(_8908_), .Y(_8924_) );
	NAND3X1 NAND3X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8924_), .C(divider_divuResult_3_bF_buf7), .Y(_8925_) );
	NAND2X1 NAND2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8496_), .Y(_8926_) );
	INVX1 INVX1_1276 ( .gnd(gnd), .vdd(vdd), .A(_8926_), .Y(_8928_) );
	NAND2X1 NAND2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .B(_8664__bF_buf6), .Y(_8929_) );
	NAND3X1 NAND3X1_1930 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf4), .B(_8929_), .C(_8925_), .Y(_8930_) );
	NAND2X1 NAND2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_8930_), .B(_8923_), .Y(_8931_) );
	NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_8919_), .Y(_8932_) );
	OAI21X1 OAI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_8516_), .B(_8517_), .C(_8664__bF_buf5), .Y(_8933_) );
	NAND2X1 NAND2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_8518_), .B(_8515_), .Y(_8934_) );
	INVX1 INVX1_1277 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .Y(_8935_) );
	AOI21X1 AOI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_8523_), .B(_8526_), .C(_8282_), .Y(_8936_) );
	OAI21X1 OAI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_8935_), .B(_8936_), .C(_8934_), .Y(_8937_) );
	INVX1 INVX1_1278 ( .gnd(gnd), .vdd(vdd), .A(_8934_), .Y(_8939_) );
	NAND2X1 NAND2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_8526_), .B(_8523_), .Y(_8940_) );
	OAI21X1 OAI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_8281_), .B(_8692_), .C(_8940_), .Y(_8941_) );
	NAND3X1 NAND3X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_8939_), .B(_8539_), .C(_8941_), .Y(_8942_) );
	NAND2X1 NAND2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_8937_), .Y(_8943_) );
	NAND2X1 NAND2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf6), .B(_8943_), .Y(_8944_) );
	NAND3X1 NAND3X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf0), .B(_8933_), .C(_8944_), .Y(_8945_) );
	NAND2X1 NAND2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_8664__bF_buf4), .Y(_8946_) );
	NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_8940_), .B(_8636_), .Y(_8947_) );
	NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(_8947_), .Y(_8948_) );
	NAND2X1 NAND2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_8948_), .B(divider_divuResult_3_bF_buf5), .Y(_8950_) );
	NAND2X1 NAND2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_8946_), .Y(_8951_) );
	NAND2X1 NAND2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf2), .B(_8951_), .Y(_8952_) );
	AOI21X1 AOI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8933_), .C(_1944__bF_buf4), .Y(_8953_) );
	OAI21X1 OAI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_8953_), .B(_8952_), .C(_8945_), .Y(_8954_) );
	OAI21X1 OAI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_8919_), .C(_8912_), .Y(_8955_) );
	AOI21X1 AOI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_8932_), .B(_8954_), .C(_8955_), .Y(_8956_) );
	NAND3X1 NAND3X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf2), .B(_8870_), .C(_8877_), .Y(_8957_) );
	AOI21X1 AOI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_8877_), .B(_8870_), .C(_3789__bF_buf1), .Y(_8958_) );
	OAI21X1 OAI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_8664__bF_buf3), .B(_8887_), .C(_8892_), .Y(_8959_) );
	NAND2X1 NAND2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf3), .B(_8959_), .Y(_8961_) );
	OAI21X1 OAI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_8961_), .B(_8958_), .C(_8957_), .Y(_8962_) );
	NAND3X1 NAND3X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf2), .B(_8834_), .C(_8847_), .Y(_8963_) );
	AOI21X1 AOI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .B(_8834_), .C(_4424__bF_buf1), .Y(_8964_) );
	AOI21X1 AOI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_8865_), .B(_8866_), .C(divider_absoluteValue_B_flipSign_result_20_bF_buf0), .Y(_8965_) );
	INVX1 INVX1_1279 ( .gnd(gnd), .vdd(vdd), .A(_8965_), .Y(_8966_) );
	OAI21X1 OAI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(_8964_), .C(_8963_), .Y(_8967_) );
	AOI21X1 AOI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .B(_8962_), .C(_8967_), .Y(_8968_) );
	OAI21X1 OAI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_8896_), .B(_8956_), .C(_8968_), .Y(_8969_) );
	AOI21X1 AOI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_8832_), .B(_8969_), .C(_8815_), .Y(_8970_) );
	OAI21X1 OAI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_8052__bF_buf0), .B(_8056_), .C(_8053_), .Y(_8972_) );
	NAND2X1 NAND2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_8972_), .B(_8664__bF_buf2), .Y(_8973_) );
	NAND2X1 NAND2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_8072_), .B(_8073_), .Y(_8974_) );
	NAND2X1 NAND2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_8076_), .B(_8079_), .Y(_8975_) );
	INVX1 INVX1_1280 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .Y(_8976_) );
	INVX1 INVX1_1281 ( .gnd(gnd), .vdd(vdd), .A(_8604_), .Y(_8977_) );
	NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_8976_), .B(_8977_), .Y(_8978_) );
	OAI21X1 OAI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_8069_), .B(_8978_), .C(_8974_), .Y(_8979_) );
	NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_8069_), .B(_8978_), .Y(_8980_) );
	OAI21X1 OAI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_8055_), .B(_8595_), .C(_8980_), .Y(_8981_) );
	NAND2X1 NAND2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_8979_), .B(_8981_), .Y(_8983_) );
	NAND2X1 NAND2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_8983_), .B(divider_divuResult_3_bF_buf4), .Y(_8984_) );
	NAND3X1 NAND3X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf6), .B(_8984_), .C(_8973_), .Y(_8985_) );
	INVX1 INVX1_1282 ( .gnd(gnd), .vdd(vdd), .A(_8978_), .Y(_8986_) );
	NAND2X1 NAND2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_8976_), .B(_8977_), .Y(_8987_) );
	NAND2X1 NAND2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_8987_), .B(_8986_), .Y(_8988_) );
	NAND2X1 NAND2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_8988_), .B(divider_divuResult_3_bF_buf3), .Y(_8989_) );
	NAND2X1 NAND2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_8068_), .B(_8664__bF_buf1), .Y(_8990_) );
	NAND3X1 NAND3X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf5), .B(_8989_), .C(_8990_), .Y(_8991_) );
	AOI21X1 AOI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_8973_), .B(_8984_), .C(_4100__bF_buf5), .Y(_8992_) );
	OAI21X1 OAI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(_8992_), .C(_8985_), .Y(_8994_) );
	INVX1 INVX1_1283 ( .gnd(gnd), .vdd(vdd), .A(_8994_), .Y(_8995_) );
	AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_8107_), .B(_8110_), .Y(_8996_) );
	INVX1 INVX1_1284 ( .gnd(gnd), .vdd(vdd), .A(_8602_), .Y(_8997_) );
	OAI21X1 OAI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf5), .B(_8997_), .C(_8601_), .Y(_8998_) );
	XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_8996_), .Y(_8999_) );
	NAND3X1 NAND3X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_8999_), .C(_8659_), .Y(_9000_) );
	OAI21X1 OAI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(divider_divuResult_3_bF_buf2), .C(_9000_), .Y(_9001_) );
	INVX1 INVX1_1285 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .Y(_9002_) );
	NAND2X1 NAND2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_8099_), .B(_8106_), .Y(_9003_) );
	XNOR2X1 XNOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_9003_), .B(_8097_), .Y(_9005_) );
	INVX1 INVX1_1286 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .Y(_9006_) );
	NAND2X1 NAND2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_9006_), .B(divider_divuResult_3_bF_buf1), .Y(_9007_) );
	NAND2X1 NAND2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(_8664__bF_buf0), .Y(_9008_) );
	NAND3X1 NAND3X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf7), .B(_9007_), .C(_9008_), .Y(_9009_) );
	OAI21X1 OAI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf6), .B(_9001_), .C(_9009_), .Y(_9010_) );
	OAI21X1 OAI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf7), .B(_9002_), .C(_9010_), .Y(_9011_) );
	INVX1 INVX1_1287 ( .gnd(gnd), .vdd(vdd), .A(_8972_), .Y(_9012_) );
	NAND2X1 NAND2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_9012_), .B(_8664__bF_buf6), .Y(_9013_) );
	INVX1 INVX1_1288 ( .gnd(gnd), .vdd(vdd), .A(_8983_), .Y(_9014_) );
	NAND2X1 NAND2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_9014_), .B(divider_divuResult_3_bF_buf0), .Y(_9016_) );
	AOI21X1 AOI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_9013_), .B(_9016_), .C(_4100__bF_buf4), .Y(_9017_) );
	AOI21X1 AOI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_8973_), .B(_8984_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf5), .Y(_9018_) );
	INVX1 INVX1_1289 ( .gnd(gnd), .vdd(vdd), .A(_8988_), .Y(_9019_) );
	NAND2X1 NAND2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_9019_), .B(divider_divuResult_3_bF_buf7), .Y(_9020_) );
	NAND2X1 NAND2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_8596_), .B(_8664__bF_buf5), .Y(_9021_) );
	AOI21X1 AOI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_9021_), .B(_9020_), .C(_1735__bF_buf4), .Y(_9022_) );
	AOI21X1 AOI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_8990_), .B(_8989_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf3), .Y(_9023_) );
	OAI22X1 OAI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_9017_), .B(_9018_), .C(_9022_), .D(_9023_), .Y(_9024_) );
	OAI21X1 OAI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_9024_), .B(_9011_), .C(_8995_), .Y(_9025_) );
	AOI21X1 AOI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_8586_), .B(_8660_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf4), .Y(_9027_) );
	NAND3X1 NAND3X1_1939 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf3), .B(_8660_), .C(_8586_), .Y(_9028_) );
	NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_2_), .B(_1746__bF_buf3), .Y(_9029_) );
	INVX1 INVX1_1290 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .Y(_9030_) );
	AOI21X1 AOI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_9028_), .B(_9030_), .C(_9027_), .Y(_9031_) );
	NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf6), .B(_9001_), .Y(_9032_) );
	INVX1 INVX1_1291 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .Y(_9033_) );
	NAND2X1 NAND2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_9033_), .B(_8664__bF_buf4), .Y(_9034_) );
	AOI21X1 AOI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_9000_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf5), .Y(_9035_) );
	NAND2X1 NAND2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(divider_divuResult_3_bF_buf6), .Y(_9036_) );
	NAND2X1 NAND2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_8602_), .B(_8664__bF_buf3), .Y(_9038_) );
	AOI21X1 AOI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_9038_), .B(_9036_), .C(_2547__bF_buf6), .Y(_9039_) );
	AOI21X1 AOI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_9008_), .B(_9007_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf6), .Y(_9040_) );
	OAI22X1 OAI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_9039_), .B(_9040_), .C(_9035_), .D(_9032_), .Y(_9041_) );
	NOR3X1 NOR3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_9024_), .C(_9041_), .Y(_9042_) );
	OAI21X1 OAI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_8153_), .B(_8156_), .C(_8664__bF_buf2), .Y(_9043_) );
	NAND2X1 NAND2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_8152_), .B(_8157_), .Y(_9044_) );
	INVX1 INVX1_1292 ( .gnd(gnd), .vdd(vdd), .A(_8200_), .Y(_9045_) );
	NAND2X1 NAND2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_8607_), .B(_8113_), .Y(_9046_) );
	AOI21X1 AOI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_9046_), .B(_8279_), .C(_9045_), .Y(_9047_) );
	OAI21X1 OAI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_8267_), .B(_9047_), .C(_8611_), .Y(_9049_) );
	NAND3X1 NAND3X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_9044_), .B(_8262_), .C(_9049_), .Y(_9050_) );
	INVX1 INVX1_1293 ( .gnd(gnd), .vdd(vdd), .A(_9044_), .Y(_9051_) );
	INVX1 INVX1_1294 ( .gnd(gnd), .vdd(vdd), .A(_8611_), .Y(_9052_) );
	AOI21X1 AOI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_8691_), .B(_8112_), .C(_8254_), .Y(_9053_) );
	OAI21X1 OAI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_8634_), .B(_9053_), .C(_8200_), .Y(_9054_) );
	AOI21X1 AOI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_9054_), .B(_8620_), .C(_9052_), .Y(_9055_) );
	OAI21X1 OAI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(_9055_), .C(_9051_), .Y(_9056_) );
	NAND3X1 NAND3X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_9056_), .B(divider_divuResult_3_bF_buf5), .C(_9050_), .Y(_9057_) );
	NAND3X1 NAND3X1_1942 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_9043_), .C(_9057_), .Y(_9058_) );
	OAI21X1 OAI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_8150_), .B(_8151_), .C(_8664__bF_buf1), .Y(_9060_) );
	OAI21X1 OAI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_8614_), .B(_9055_), .C(_9044_), .Y(_9061_) );
	NAND3X1 NAND3X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_9051_), .B(_8262_), .C(_9049_), .Y(_9062_) );
	NAND3X1 NAND3X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(divider_divuResult_3_bF_buf4), .C(_9062_), .Y(_9063_) );
	NAND3X1 NAND3X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf0), .B(_9060_), .C(_9063_), .Y(_9064_) );
	INVX1 INVX1_1295 ( .gnd(gnd), .vdd(vdd), .A(_8264_), .Y(_9065_) );
	OAI21X1 OAI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_8254_), .B(_8605_), .C(_8279_), .Y(_9066_) );
	AOI22X1 AOI22X1_199 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_8619_), .C(_8200_), .D(_9066_), .Y(_9067_) );
	NAND2X1 NAND2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_9052_), .B(_9067_), .Y(_9068_) );
	NAND2X1 NAND2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_9068_), .B(_9049_), .Y(_9069_) );
	NAND2X1 NAND2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_9069_), .B(divider_divuResult_3_bF_buf3), .Y(_9071_) );
	INVX1 INVX1_1296 ( .gnd(gnd), .vdd(vdd), .A(_8261_), .Y(_9072_) );
	NAND2X1 NAND2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_9072_), .B(_8664__bF_buf0), .Y(_9073_) );
	NAND3X1 NAND3X1_1946 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .B(_9071_), .C(_9073_), .Y(_9074_) );
	XNOR2X1 XNOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_9067_), .B(_8611_), .Y(_9075_) );
	NAND2X1 NAND2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf2), .B(_9075_), .Y(_9076_) );
	NAND2X1 NAND2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_8261_), .B(_8664__bF_buf6), .Y(_9077_) );
	NAND3X1 NAND3X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf2), .B(_9077_), .C(_9076_), .Y(_9078_) );
	AOI22X1 AOI22X1_200 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_9074_), .C(_9058_), .D(_9064_), .Y(_9079_) );
	NAND2X1 NAND2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .B(_8664__bF_buf5), .Y(_9080_) );
	NAND2X1 NAND2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_8180_), .B(_8186_), .Y(_9082_) );
	INVX1 INVX1_1297 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .Y(_9083_) );
	AOI22X1 AOI22X1_201 ( .gnd(gnd), .vdd(vdd), .A(_8195_), .B(_8199_), .C(_8279_), .D(_9046_), .Y(_9084_) );
	OAI21X1 OAI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_9083_), .B(_9084_), .C(_9082_), .Y(_9085_) );
	INVX1 INVX1_1298 ( .gnd(gnd), .vdd(vdd), .A(_9082_), .Y(_9086_) );
	NAND2X1 NAND2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_8199_), .B(_8195_), .Y(_9087_) );
	OAI21X1 OAI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_8634_), .B(_9053_), .C(_9087_), .Y(_9088_) );
	NAND3X1 NAND3X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_9086_), .B(_8266_), .C(_9088_), .Y(_9089_) );
	NAND2X1 NAND2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_9085_), .Y(_9090_) );
	NAND2X1 NAND2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_9090_), .B(divider_divuResult_3_bF_buf1), .Y(_9091_) );
	NAND3X1 NAND3X1_1949 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf1), .B(_9091_), .C(_9080_), .Y(_9093_) );
	NAND2X1 NAND2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .B(_8664__bF_buf4), .Y(_9094_) );
	NAND3X1 NAND3X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_9085_), .B(_9089_), .C(divider_divuResult_3_bF_buf0), .Y(_9095_) );
	NAND3X1 NAND3X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf1), .B(_9094_), .C(_9095_), .Y(_9096_) );
	NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_9066_), .Y(_9097_) );
	NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(_9097_), .Y(_9098_) );
	INVX1 INVX1_1299 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .Y(_9099_) );
	NAND2X1 NAND2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_9099_), .B(divider_divuResult_3_bF_buf7), .Y(_9100_) );
	NAND2X1 NAND2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .B(_8664__bF_buf3), .Y(_9101_) );
	NAND3X1 NAND3X1_1952 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .B(_9100_), .C(_9101_), .Y(_9102_) );
	NAND3X1 NAND3X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_9098_), .C(_8659_), .Y(_9104_) );
	INVX1 INVX1_1300 ( .gnd(gnd), .vdd(vdd), .A(_8618_), .Y(_9105_) );
	NAND2X1 NAND2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .B(_8664__bF_buf2), .Y(_9106_) );
	NAND3X1 NAND3X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf3), .B(_9104_), .C(_9106_), .Y(_9107_) );
	AOI22X1 AOI22X1_202 ( .gnd(gnd), .vdd(vdd), .A(_9102_), .B(_9107_), .C(_9093_), .D(_9096_), .Y(_9108_) );
	NAND2X1 NAND2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_9079_), .Y(_9109_) );
	OAI21X1 OAI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_8212_), .B(_8213_), .C(_8664__bF_buf1), .Y(_9110_) );
	NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf6), .B(_8273_), .Y(_9111_) );
	INVX1 INVX1_1301 ( .gnd(gnd), .vdd(vdd), .A(_8228_), .Y(_9112_) );
	NAND2X1 NAND2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_8253_), .B(_8113_), .Y(_9113_) );
	AOI21X1 AOI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_9113_), .B(_8633_), .C(_9112_), .Y(_9115_) );
	OAI21X1 OAI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_9111_), .B(_9115_), .C(_8216_), .Y(_9116_) );
	INVX1 INVX1_1302 ( .gnd(gnd), .vdd(vdd), .A(_8216_), .Y(_9117_) );
	INVX1 INVX1_1303 ( .gnd(gnd), .vdd(vdd), .A(_9111_), .Y(_9118_) );
	NAND2X1 NAND2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_8633_), .B(_9113_), .Y(_9119_) );
	NAND2X1 NAND2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_8228_), .B(_9119_), .Y(_9120_) );
	NAND3X1 NAND3X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(_9118_), .C(_9120_), .Y(_9121_) );
	NAND2X1 NAND2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_9116_), .B(_9121_), .Y(_9122_) );
	NAND2X1 NAND2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf6), .B(_9122_), .Y(_9123_) );
	NAND3X1 NAND3X1_1956 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf0), .B(_9110_), .C(_9123_), .Y(_9124_) );
	AOI21X1 AOI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_8659_), .B(_2020_), .C(_8626_), .Y(_9126_) );
	AOI21X1 AOI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_9116_), .B(_9121_), .C(_8664__bF_buf0), .Y(_9127_) );
	OAI21X1 OAI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_9127_), .C(_8971__bF_buf5), .Y(_9128_) );
	NAND2X1 NAND2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_9124_), .B(_9128_), .Y(_9129_) );
	NAND3X1 NAND3X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8633_), .C(_9113_), .Y(_9130_) );
	NAND2X1 NAND2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_9130_), .B(_9120_), .Y(_9131_) );
	NAND2X1 NAND2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_9131_), .B(divider_divuResult_3_bF_buf5), .Y(_9132_) );
	NAND2X1 NAND2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_8273_), .B(_8664__bF_buf6), .Y(_9133_) );
	NAND3X1 NAND3X1_1958 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .B(_9132_), .C(_9133_), .Y(_9134_) );
	INVX1 INVX1_1304 ( .gnd(gnd), .vdd(vdd), .A(_9131_), .Y(_9135_) );
	NAND2X1 NAND2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_9135_), .B(divider_divuResult_3_bF_buf4), .Y(_9137_) );
	INVX1 INVX1_1305 ( .gnd(gnd), .vdd(vdd), .A(_8273_), .Y(_9138_) );
	NAND2X1 NAND2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_9138_), .B(_8664__bF_buf5), .Y(_9139_) );
	NAND3X1 NAND3X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf2), .B(_9137_), .C(_9139_), .Y(_9140_) );
	NAND2X1 NAND2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_9134_), .B(_9140_), .Y(_9141_) );
	NAND2X1 NAND2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_8252_), .B(_8249_), .Y(_9142_) );
	XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_8113_), .B(_9142_), .Y(_9143_) );
	INVX1 INVX1_1306 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .Y(_9144_) );
	NAND3X1 NAND3X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_9144_), .C(_8659_), .Y(_9145_) );
	NAND2X1 NAND2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_8630_), .B(_8664__bF_buf4), .Y(_9146_) );
	NAND3X1 NAND3X1_1961 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .B(_9145_), .C(_9146_), .Y(_9148_) );
	INVX1 INVX1_1307 ( .gnd(gnd), .vdd(vdd), .A(_8630_), .Y(_9149_) );
	NAND2X1 NAND2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .B(_8664__bF_buf3), .Y(_9150_) );
	NAND3X1 NAND3X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_9143_), .C(_8659_), .Y(_9151_) );
	NAND3X1 NAND3X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf5), .B(_9151_), .C(_9150_), .Y(_9152_) );
	NAND2X1 NAND2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_8628_), .B(_8664__bF_buf2), .Y(_9153_) );
	NAND2X1 NAND2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_8238_), .B(_8243_), .Y(_9154_) );
	NAND2X1 NAND2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_9142_), .B(_8113_), .Y(_9155_) );
	AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_9155_), .B(_8277_), .Y(_9156_) );
	AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_9156_), .B(_9154_), .Y(_9157_) );
	NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_9156_), .Y(_9159_) );
	NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_9159_), .B(_9157_), .Y(_9160_) );
	NAND2X1 NAND2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf3), .B(_9160_), .Y(_9161_) );
	NAND3X1 NAND3X1_1964 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf5), .B(_9153_), .C(_9161_), .Y(_9162_) );
	NAND3X1 NAND3X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_8229_), .B(_8237_), .C(_8664__bF_buf1), .Y(_9163_) );
	OAI21X1 OAI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_9157_), .B(_9159_), .C(divider_divuResult_3_bF_buf2), .Y(_9164_) );
	NAND3X1 NAND3X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf4), .B(_9164_), .C(_9163_), .Y(_9165_) );
	AOI22X1 AOI22X1_203 ( .gnd(gnd), .vdd(vdd), .A(_9148_), .B(_9152_), .C(_9162_), .D(_9165_), .Y(_9166_) );
	NAND3X1 NAND3X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_9141_), .B(_9129_), .C(_9166_), .Y(_9167_) );
	NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_9109_), .B(_9167_), .Y(_9168_) );
	OAI21X1 OAI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_9025_), .B(_9042_), .C(_9168_), .Y(_9170_) );
	AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_9079_), .B(_9108_), .Y(_9171_) );
	NOR3X1 NOR3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf4), .B(_9126_), .C(_9127_), .Y(_9172_) );
	AOI21X1 AOI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_9110_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf6), .Y(_9173_) );
	OAI21X1 OAI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_9172_), .B(_9173_), .C(_9141_), .Y(_9174_) );
	NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_9127_), .Y(_9175_) );
	NAND3X1 NAND3X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf3), .B(_9110_), .C(_9123_), .Y(_9176_) );
	OAI21X1 OAI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_9138_), .B(divider_divuResult_3_bF_buf1), .C(_9132_), .Y(_9177_) );
	OAI21X1 OAI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_9177_), .C(_9176_), .Y(_9178_) );
	OAI21X1 OAI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf2), .B(_9175_), .C(_9178_), .Y(_9179_) );
	AOI21X1 AOI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_9150_), .B(_9151_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .Y(_9181_) );
	AOI21X1 AOI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_9163_), .B(_9164_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf4), .Y(_9182_) );
	NAND3X1 NAND3X1_1969 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf3), .B(_9164_), .C(_9163_), .Y(_9183_) );
	OAI21X1 OAI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_9181_), .B(_9182_), .C(_9183_), .Y(_9184_) );
	OAI21X1 OAI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_9184_), .B(_9174_), .C(_9179_), .Y(_9185_) );
	NAND2X1 NAND2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(_9064_), .Y(_9186_) );
	NAND2X1 NAND2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_9074_), .B(_9078_), .Y(_9187_) );
	NAND2X1 NAND2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .B(_9186_), .Y(_9188_) );
	OAI21X1 OAI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_8664__bF_buf0), .B(_9090_), .C(_9094_), .Y(_9189_) );
	OAI21X1 OAI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_8617_), .B(divider_divuResult_3_bF_buf0), .C(_9091_), .Y(_9190_) );
	NAND3X1 NAND3X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf2), .B(_9100_), .C(_9101_), .Y(_9192_) );
	OAI21X1 OAI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf0), .B(_9190_), .C(_9192_), .Y(_9193_) );
	OAI21X1 OAI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf0), .B(_9189_), .C(_9193_), .Y(_9194_) );
	AOI21X1 AOI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_9063_), .B(_9060_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .Y(_9195_) );
	NAND3X1 NAND3X1_1971 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf3), .B(_9060_), .C(_9063_), .Y(_9196_) );
	AOI21X1 AOI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_9076_), .B(_9077_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf4), .Y(_9197_) );
	AOI21X1 AOI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_9196_), .C(_9195_), .Y(_9198_) );
	OAI21X1 OAI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_9194_), .C(_9198_), .Y(_9199_) );
	AOI21X1 AOI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_9171_), .C(_9199_), .Y(_9200_) );
	NAND2X1 NAND2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_9200_), .B(_9170_), .Y(_9201_) );
	NAND3X1 NAND3X1_1972 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf2), .B(_8851_), .C(_8854_), .Y(_9203_) );
	NAND2X1 NAND2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_8867_), .B(_8863_), .Y(_9204_) );
	NAND3X1 NAND3X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_8963_), .B(_9203_), .C(_9204_), .Y(_9205_) );
	NAND3X1 NAND3X1_1974 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf0), .B(_8880_), .C(_8884_), .Y(_9206_) );
	NAND2X1 NAND2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_8893_), .B(_8890_), .Y(_9207_) );
	NAND3X1 NAND3X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_9207_), .B(_9206_), .C(_8957_), .Y(_9208_) );
	NAND3X1 NAND3X1_1976 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf4), .B(_8897_), .C(_8911_), .Y(_9209_) );
	NAND3X1 NAND3X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf3), .B(_8913_), .C(_8917_), .Y(_9210_) );
	NAND2X1 NAND2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_9209_), .B(_9210_), .Y(_9211_) );
	AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_8930_), .Y(_9212_) );
	NAND3X1 NAND3X1_1978 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf4), .B(_8933_), .C(_8944_), .Y(_9214_) );
	NAND2X1 NAND2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_8514_), .B(_8513_), .Y(_9215_) );
	INVX1 INVX1_1308 ( .gnd(gnd), .vdd(vdd), .A(_9215_), .Y(_9216_) );
	NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_9216_), .B(divider_divuResult_3_bF_buf7), .Y(_9217_) );
	AOI21X1 AOI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_8937_), .B(_8942_), .C(_8664__bF_buf6), .Y(_9218_) );
	OAI21X1 OAI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(_9218_), .C(_1944__bF_buf3), .Y(_9219_) );
	OAI21X1 OAI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(_8947_), .C(divider_divuResult_3_bF_buf6), .Y(_9220_) );
	NAND3X1 NAND3X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_8524_), .B(_8525_), .C(_8664__bF_buf5), .Y(_9221_) );
	NAND3X1 NAND3X1_1980 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf1), .B(_9220_), .C(_9221_), .Y(_9222_) );
	NAND3X1 NAND3X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf1), .B(_8950_), .C(_8946_), .Y(_9223_) );
	AOI22X1 AOI22X1_204 ( .gnd(gnd), .vdd(vdd), .A(_9222_), .B(_9223_), .C(_9214_), .D(_9219_), .Y(_9225_) );
	NAND3X1 NAND3X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_9212_), .B(_9211_), .C(_9225_), .Y(_9226_) );
	NOR3X1 NOR3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_9226_), .C(_9205_), .Y(_9227_) );
	NAND3X1 NAND3X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_9227_), .B(_8832_), .C(_9201_), .Y(_9228_) );
	AOI21X1 AOI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_8970_), .B(_9228_), .C(_8663_), .Y(divider_divuResult_2_) );
	NAND2X1 NAND2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_3_), .B(_1746__bF_buf2), .Y(_9229_) );
	NAND3X1 NAND3X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_9229_), .C(divider_divuResult_3_bF_buf5), .Y(_9230_) );
	NAND2X1 NAND2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_8587_), .B(_8664__bF_buf4), .Y(_9231_) );
	AOI21X1 AOI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_9230_), .B(_9231_), .C(_1768__bF_buf6), .Y(_9232_) );
	NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_9027_), .B(_9232_), .Y(_9233_) );
	XNOR2X1 XNOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_9233_), .B(_9029_), .Y(_9235_) );
	INVX1 INVX1_1309 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .Y(_9236_) );
	NAND2X1 NAND2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_9236_), .B(divider_divuResult_2_bF_buf7), .Y(_9237_) );
	OAI21X1 OAI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_8661_), .B(divider_divuResult_2_bF_buf6), .C(_9237_), .Y(_9238_) );
	NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf5), .B(_9238_), .Y(_9239_) );
	INVX1 INVX1_1310 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .Y(_9240_) );
	NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_8819_), .B(_8822_), .Y(_9241_) );
	NAND3X1 NAND3X1_1985 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_8757_), .C(_8760_), .Y(_9242_) );
	NAND2X1 NAND2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_8774_), .B(_8768_), .Y(_9243_) );
	NAND3X1 NAND3X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_8799_), .B(_9242_), .C(_9243_), .Y(_9244_) );
	NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_8777_), .B(_8789_), .Y(_9246_) );
	OAI21X1 OAI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf1), .B(_9246_), .C(_8797_), .Y(_9247_) );
	INVX1 INVX1_1311 ( .gnd(gnd), .vdd(vdd), .A(_8799_), .Y(_9248_) );
	INVX1 INVX1_1312 ( .gnd(gnd), .vdd(vdd), .A(_8801_), .Y(_9249_) );
	AOI21X1 AOI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_9249_), .B(_9242_), .C(_9248_), .Y(_9250_) );
	OAI21X1 OAI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_9244_), .B(_9247_), .C(_9250_), .Y(_9251_) );
	NOR3X1 NOR3X1_93 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_8729_), .C(_8732_), .Y(_9252_) );
	INVX1 INVX1_1313 ( .gnd(gnd), .vdd(vdd), .A(_8807_), .Y(_9253_) );
	AOI21X1 AOI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_8820_), .B(_9253_), .C(_9252_), .Y(_9254_) );
	AOI21X1 AOI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_8714_), .B(_8715_), .C(divider_absoluteValue_B_flipSign_result_28_), .Y(_9255_) );
	AOI21X1 AOI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_8816_), .C(_8809_), .Y(_9257_) );
	OAI21X1 OAI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_8819_), .B(_9254_), .C(_9257_), .Y(_9258_) );
	AOI21X1 AOI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .B(_9241_), .C(_9258_), .Y(_9259_) );
	AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_8827_), .B(_8826_), .Y(_9260_) );
	NAND3X1 NAND3X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_8790_), .B(_8791_), .C(_9260_), .Y(_9261_) );
	NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_9244_), .B(_9261_), .Y(_9262_) );
	NAND2X1 NAND2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_9262_), .B(_9241_), .Y(_9263_) );
	NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_9205_), .Y(_9264_) );
	NAND3X1 NAND3X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_9211_), .B(_9212_), .C(_8954_), .Y(_9265_) );
	OAI21X1 OAI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_8543_), .B(divider_divuResult_3_bF_buf4), .C(_8911_), .Y(_9266_) );
	INVX1 INVX1_1314 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .Y(_9268_) );
	INVX1 INVX1_1315 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .Y(_9269_) );
	OAI21X1 OAI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf2), .B(_9268_), .C(_9269_), .Y(_9270_) );
	NAND3X1 NAND3X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_8912_), .B(_9270_), .C(_9265_), .Y(_9271_) );
	AOI21X1 AOI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .B(_8880_), .C(divider_absoluteValue_B_flipSign_result_19_bF_buf4), .Y(_9272_) );
	INVX1 INVX1_1316 ( .gnd(gnd), .vdd(vdd), .A(_8961_), .Y(_9273_) );
	AOI21X1 AOI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .B(_9206_), .C(_9272_), .Y(_9274_) );
	AOI21X1 AOI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8851_), .C(divider_absoluteValue_B_flipSign_result_21_bF_buf1), .Y(_9275_) );
	AOI21X1 AOI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_8965_), .B(_9203_), .C(_9275_), .Y(_9276_) );
	OAI21X1 OAI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_9274_), .B(_9205_), .C(_9276_), .Y(_9277_) );
	AOI21X1 AOI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_9264_), .B(_9271_), .C(_9277_), .Y(_9279_) );
	OAI21X1 OAI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_9263_), .B(_9279_), .C(_9259_), .Y(_9280_) );
	NAND3X1 NAND3X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf5), .B(_9000_), .C(_9034_), .Y(_9281_) );
	AOI21X1 AOI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_9000_), .C(_2470__bF_buf4), .Y(_9282_) );
	OAI21X1 OAI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_9009_), .B(_9282_), .C(_9281_), .Y(_9283_) );
	NAND3X1 NAND3X1_1991 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf4), .B(_8984_), .C(_8973_), .Y(_9284_) );
	NAND3X1 NAND3X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf3), .B(_9016_), .C(_9013_), .Y(_9285_) );
	NAND3X1 NAND3X1_1993 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf2), .B(_8989_), .C(_8990_), .Y(_9286_) );
	NAND3X1 NAND3X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_9020_), .C(_9021_), .Y(_9287_) );
	AOI22X1 AOI22X1_205 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9285_), .C(_9286_), .D(_9287_), .Y(_9288_) );
	AOI21X1 AOI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_9283_), .B(_9288_), .C(_8994_), .Y(_9290_) );
	NAND2X1 NAND2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf5), .B(_8661_), .Y(_9291_) );
	OAI21X1 OAI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_9232_), .C(_9291_), .Y(_9292_) );
	NAND3X1 NAND3X1_1995 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf4), .B(_9000_), .C(_9034_), .Y(_9293_) );
	NAND2X1 NAND2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf3), .B(_9001_), .Y(_9294_) );
	NAND3X1 NAND3X1_1996 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf4), .B(_9007_), .C(_9008_), .Y(_9295_) );
	NAND3X1 NAND3X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf5), .B(_9036_), .C(_9038_), .Y(_9296_) );
	AOI22X1 AOI22X1_206 ( .gnd(gnd), .vdd(vdd), .A(_9296_), .B(_9295_), .C(_9293_), .D(_9294_), .Y(_9297_) );
	NAND3X1 NAND3X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .B(_9297_), .C(_9292_), .Y(_9298_) );
	NAND2X1 NAND2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .B(_9290_), .Y(_9299_) );
	OAI21X1 OAI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_9127_), .C(divider_absoluteValue_B_flipSign_result_9_bF_buf5), .Y(_9301_) );
	AOI22X1 AOI22X1_207 ( .gnd(gnd), .vdd(vdd), .A(_9134_), .B(_9140_), .C(_9124_), .D(_9128_), .Y(_9302_) );
	OAI21X1 OAI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_8630_), .B(divider_divuResult_3_bF_buf3), .C(_9151_), .Y(_9303_) );
	NAND2X1 NAND2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf4), .B(_9303_), .Y(_9304_) );
	NAND3X1 NAND3X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf3), .B(_9153_), .C(_9161_), .Y(_9305_) );
	AOI21X1 AOI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_9153_), .C(_4714__bF_buf2), .Y(_9306_) );
	AOI21X1 AOI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_9305_), .C(_9306_), .Y(_9307_) );
	AOI22X1 AOI22X1_208 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .B(_9178_), .C(_9307_), .D(_9302_), .Y(_9308_) );
	NAND3X1 NAND3X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf5), .B(_9091_), .C(_9080_), .Y(_9309_) );
	AOI21X1 AOI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_9080_), .B(_9091_), .C(_1265__bF_buf4), .Y(_9310_) );
	OAI21X1 OAI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_9192_), .B(_9310_), .C(_9309_), .Y(_9312_) );
	OAI21X1 OAI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_8260_), .B(divider_divuResult_3_bF_buf2), .C(_9063_), .Y(_9313_) );
	NAND2X1 NAND2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf4), .B(_9313_), .Y(_9314_) );
	AOI21X1 AOI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_9057_), .B(_9043_), .C(_1494__bF_buf3), .Y(_9315_) );
	OAI21X1 OAI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_8664__bF_buf3), .B(_9069_), .C(_9077_), .Y(_9316_) );
	NAND2X1 NAND2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf1), .B(_9316_), .Y(_9317_) );
	OAI21X1 OAI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .B(_9317_), .C(_9314_), .Y(_9318_) );
	AOI21X1 AOI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .B(_9079_), .C(_9318_), .Y(_9319_) );
	OAI21X1 OAI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_9109_), .B(_9308_), .C(_9319_), .Y(_9320_) );
	AOI21X1 AOI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9168_), .C(_9320_), .Y(_9321_) );
	NAND3X1 NAND3X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_9262_), .B(_9241_), .C(_9227_), .Y(_9323_) );
	NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_9323_), .Y(_9324_) );
	OAI21X1 OAI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .B(_9280_), .C(_8662_), .Y(_9325_) );
	NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .B(_9325__bF_buf6), .Y(_9326_) );
	NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_8661_), .B(divider_divuResult_2_bF_buf5), .Y(_9327_) );
	OAI21X1 OAI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9326_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf3), .Y(_9328_) );
	INVX1 INVX1_1317 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .Y(_9329_) );
	OAI21X1 OAI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_1746__bF_buf1), .B(_9325__bF_buf5), .C(divider_aOp_abs_2_), .Y(_9330_) );
	NAND2X1 NAND2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(divider_divuResult_2_bF_buf4), .Y(_9331_) );
	AOI21X1 AOI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_9330_), .B(_9331_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf2), .Y(_9332_) );
	NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_1_), .B(_1746__bF_buf0), .Y(_9334_) );
	INVX1 INVX1_1318 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .Y(_9335_) );
	NAND3X1 NAND3X1_2002 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf1), .B(_9331_), .C(_9330_), .Y(_9336_) );
	AOI21X1 AOI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .B(_9336_), .C(_9332_), .Y(_9337_) );
	OAI21X1 OAI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_9329_), .B(_9337_), .C(_9240_), .Y(_9338_) );
	NAND3X1 NAND3X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_9013_), .B(_9016_), .C(_9325__bF_buf4), .Y(_9339_) );
	NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_9022_), .B(_9023_), .Y(_9340_) );
	AOI21X1 AOI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(_9297_), .C(_9283_), .Y(_9341_) );
	OAI21X1 OAI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_9340_), .B(_9341_), .C(_8991_), .Y(_9342_) );
	OAI21X1 OAI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_9017_), .B(_9018_), .C(_9342_), .Y(_9343_) );
	NAND2X1 NAND2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_9284_), .B(_9285_), .Y(_9345_) );
	OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_9342_), .B(_9345_), .Y(_9346_) );
	NAND2X1 NAND2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_9346_), .Y(_9347_) );
	NAND2X1 NAND2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_9347_), .B(divider_divuResult_2_bF_buf3), .Y(_9348_) );
	NAND3X1 NAND3X1_2004 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf6), .B(_9348_), .C(_9339_), .Y(_9349_) );
	NAND3X1 NAND3X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_8973_), .B(_8984_), .C(_9325__bF_buf3), .Y(_9350_) );
	INVX1 INVX1_1319 ( .gnd(gnd), .vdd(vdd), .A(_9347_), .Y(_9351_) );
	NAND2X1 NAND2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_9351_), .B(divider_divuResult_2_bF_buf2), .Y(_9352_) );
	NAND3X1 NAND3X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf3), .B(_9352_), .C(_9350_), .Y(_9353_) );
	XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_9341_), .B(_9340_), .Y(_9354_) );
	INVX1 INVX1_1320 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .Y(_9356_) );
	NAND2X1 NAND2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_9356_), .B(divider_divuResult_2_bF_buf1), .Y(_9357_) );
	NAND3X1 NAND3X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .B(_9021_), .C(_9325__bF_buf2), .Y(_9358_) );
	NAND3X1 NAND3X1_2008 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf3), .B(_9357_), .C(_9358_), .Y(_9359_) );
	NAND2X1 NAND2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(divider_divuResult_2_bF_buf0), .Y(_9360_) );
	NAND3X1 NAND3X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_8989_), .B(_8990_), .C(_9325__bF_buf1), .Y(_9361_) );
	NAND3X1 NAND3X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf2), .B(_9360_), .C(_9361_), .Y(_9362_) );
	AOI22X1 AOI22X1_209 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_9349_), .C(_9359_), .D(_9362_), .Y(_9363_) );
	NAND2X1 NAND2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_8832_), .B(_8969_), .Y(_9364_) );
	NAND3X1 NAND3X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_9259_), .B(_9364_), .C(_9228_), .Y(_9365_) );
	OAI21X1 OAI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_9039_), .B(_9040_), .C(_9292_), .Y(_9367_) );
	NAND2X1 NAND2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_9296_), .Y(_9368_) );
	INVX1 INVX1_1321 ( .gnd(gnd), .vdd(vdd), .A(_9368_), .Y(_9369_) );
	NAND2X1 NAND2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_9369_), .Y(_9370_) );
	AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_9370_), .Y(_9371_) );
	INVX1 INVX1_1322 ( .gnd(gnd), .vdd(vdd), .A(_9371_), .Y(_9372_) );
	NAND3X1 NAND3X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_8662_), .B(_9372_), .C(_9365_), .Y(_9373_) );
	OAI21X1 OAI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(divider_divuResult_3_bF_buf1), .C(_9036_), .Y(_9374_) );
	INVX1 INVX1_1323 ( .gnd(gnd), .vdd(vdd), .A(_9374_), .Y(_9375_) );
	NAND2X1 NAND2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_9375_), .B(_9325__bF_buf0), .Y(_9376_) );
	NAND3X1 NAND3X1_2013 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf3), .B(_9373_), .C(_9376_), .Y(_9378_) );
	NAND2X1 NAND2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_9371_), .B(divider_divuResult_2_bF_buf7), .Y(_9379_) );
	NAND2X1 NAND2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_9374_), .B(_9325__bF_buf6), .Y(_9380_) );
	NAND3X1 NAND3X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf2), .B(_9379_), .C(_9380_), .Y(_9381_) );
	OAI21X1 OAI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_9369_), .C(_9009_), .Y(_9382_) );
	OAI21X1 OAI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_9032_), .B(_9035_), .C(_9382_), .Y(_9383_) );
	NAND2X1 NAND2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_9293_), .B(_9294_), .Y(_9384_) );
	OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_9382_), .B(_9384_), .Y(_9385_) );
	NAND2X1 NAND2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_9383_), .B(_9385_), .Y(_9386_) );
	NAND3X1 NAND3X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_8662_), .B(_9386_), .C(_9365_), .Y(_9387_) );
	NAND2X1 NAND2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_9325__bF_buf5), .Y(_9389_) );
	NAND3X1 NAND3X1_2016 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf1), .B(_9387_), .C(_9389_), .Y(_9390_) );
	OAI21X1 OAI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(divider_divuResult_2_bF_buf6), .C(_9387_), .Y(_9391_) );
	NAND2X1 NAND2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_9391_), .Y(_9392_) );
	AOI22X1 AOI22X1_210 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_9381_), .C(_9390_), .D(_9392_), .Y(_9393_) );
	AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_9393_), .B(_9363_), .Y(_9394_) );
	AOI21X1 AOI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_9350_), .B(_9352_), .C(_4999__bF_buf2), .Y(_9395_) );
	AOI21X1 AOI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_9339_), .B(_9348_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf5), .Y(_9396_) );
	AOI21X1 AOI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_9361_), .B(_9360_), .C(_4100__bF_buf1), .Y(_9397_) );
	AOI21X1 AOI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_9358_), .B(_9357_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf2), .Y(_9398_) );
	OAI22X1 OAI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_9395_), .C(_9397_), .D(_9398_), .Y(_9400_) );
	INVX1 INVX1_1324 ( .gnd(gnd), .vdd(vdd), .A(_9391_), .Y(_9401_) );
	OAI21X1 OAI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_9374_), .B(divider_divuResult_2_bF_buf5), .C(_9373_), .Y(_9402_) );
	OAI22X1 OAI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_3_bF_buf2), .B(_9402_), .C(divider_absoluteValue_B_flipSign_result_4_bF_buf0), .D(_9391_), .Y(_9403_) );
	OAI21X1 OAI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_9401_), .C(_9403_), .Y(_9404_) );
	AOI21X1 AOI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_9350_), .B(_9352_), .C(divider_absoluteValue_B_flipSign_result_6_bF_buf4), .Y(_9405_) );
	OAI21X1 OAI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf4), .B(_9351_), .C(_9339_), .Y(_9406_) );
	NAND2X1 NAND2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf3), .B(_9406_), .Y(_9407_) );
	AOI21X1 AOI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_9361_), .B(_9360_), .C(divider_absoluteValue_B_flipSign_result_5_bF_buf1), .Y(_9408_) );
	OAI21X1 OAI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_9405_), .B(_9408_), .C(_9407_), .Y(_9409_) );
	OAI21X1 OAI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_9400_), .B(_9404_), .C(_9409_), .Y(_9411_) );
	AOI21X1 AOI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_9338_), .B(_9394_), .C(_9411_), .Y(_9412_) );
	NAND3X1 NAND3X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_9060_), .B(_9063_), .C(_9325__bF_buf3), .Y(_9413_) );
	INVX1 INVX1_1325 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .Y(_9414_) );
	AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_9302_), .B(_9166_), .Y(_9415_) );
	OAI21X1 OAI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_9025_), .B(_9042_), .C(_9415_), .Y(_9416_) );
	AOI21X1 AOI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_9416_), .B(_9308_), .C(_9414_), .Y(_9417_) );
	OAI21X1 OAI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .B(_9417_), .C(_9187_), .Y(_9418_) );
	NAND3X1 NAND3X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .B(_9317_), .C(_9418_), .Y(_9419_) );
	INVX1 INVX1_1326 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .Y(_9420_) );
	INVX1 INVX1_1327 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .Y(_9422_) );
	AOI21X1 AOI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_9290_), .B(_9298_), .C(_9167_), .Y(_9423_) );
	OAI21X1 OAI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_9423_), .C(_9108_), .Y(_9424_) );
	AOI21X1 AOI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_9424_), .B(_9194_), .C(_9422_), .Y(_9425_) );
	OAI21X1 OAI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_9425_), .C(_9420_), .Y(_9426_) );
	NAND3X1 NAND3X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_9426_), .B(divider_divuResult_2_bF_buf4), .C(_9419_), .Y(_9427_) );
	NAND3X1 NAND3X1_2020 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf0), .B(_9413_), .C(_9427_), .Y(_9428_) );
	NAND2X1 NAND2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_9313_), .B(_9325__bF_buf2), .Y(_9429_) );
	OAI21X1 OAI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_9425_), .C(_9186_), .Y(_9430_) );
	NAND3X1 NAND3X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_9420_), .B(_9317_), .C(_9418_), .Y(_9431_) );
	NAND3X1 NAND3X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_9430_), .B(divider_divuResult_2_bF_buf3), .C(_9431_), .Y(_9433_) );
	NAND3X1 NAND3X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf0), .B(_9429_), .C(_9433_), .Y(_9434_) );
	NAND3X1 NAND3X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_9422_), .B(_9194_), .C(_9424_), .Y(_9435_) );
	NAND2X1 NAND2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_9435_), .B(_9418_), .Y(_9436_) );
	NAND2X1 NAND2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_9436_), .B(divider_divuResult_2_bF_buf2), .Y(_9437_) );
	OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf1), .B(_9316_), .Y(_9438_) );
	NAND3X1 NAND3X1_2025 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf2), .B(_9437_), .C(_9438_), .Y(_9439_) );
	OAI21X1 OAI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_9316_), .B(divider_divuResult_2_bF_buf0), .C(_9437_), .Y(_9440_) );
	NAND2X1 NAND2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf2), .B(_9440_), .Y(_9441_) );
	AOI22X1 AOI22X1_211 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .B(_9434_), .C(_9439_), .D(_9441_), .Y(_9442_) );
	NAND2X1 NAND2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_9093_), .B(_9096_), .Y(_9444_) );
	NAND2X1 NAND2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_9107_), .B(_9102_), .Y(_9445_) );
	INVX1 INVX1_1328 ( .gnd(gnd), .vdd(vdd), .A(_9445_), .Y(_9446_) );
	NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_9423_), .Y(_9447_) );
	OAI21X1 OAI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_9447_), .C(_9192_), .Y(_9448_) );
	XNOR2X1 XNOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_9448_), .B(_9444_), .Y(_9449_) );
	NAND2X1 NAND2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf7), .B(_9449_), .Y(_9450_) );
	NAND2X1 NAND2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_9190_), .B(_9325__bF_buf1), .Y(_9451_) );
	NAND3X1 NAND3X1_2026 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf3), .B(_9451_), .C(_9450_), .Y(_9452_) );
	XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_9448_), .B(_9444_), .Y(_9453_) );
	NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf0), .B(_9453_), .Y(_9455_) );
	NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_9189_), .B(divider_divuResult_2_bF_buf6), .Y(_9456_) );
	OAI21X1 OAI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_9456_), .B(_9455_), .C(_1484__bF_buf0), .Y(_9457_) );
	XNOR2X1 XNOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_9447_), .B(_9446_), .Y(_9458_) );
	NAND2X1 NAND2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_9458_), .B(divider_divuResult_2_bF_buf5), .Y(_9459_) );
	OAI21X1 OAI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .B(divider_divuResult_3_bF_buf0), .C(_9100_), .Y(_9460_) );
	NAND2X1 NAND2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_9460_), .B(_9325__bF_buf6), .Y(_9461_) );
	NAND3X1 NAND3X1_2027 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_11_bF_buf5), .B(_9459_), .C(_9461_), .Y(_9462_) );
	OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf5), .B(_9458_), .Y(_9463_) );
	OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf4), .B(_9460_), .Y(_9464_) );
	NAND3X1 NAND3X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf3), .B(_9464_), .C(_9463_), .Y(_9466_) );
	AOI22X1 AOI22X1_212 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_9462_), .C(_9452_), .D(_9457_), .Y(_9467_) );
	AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_9467_), .B(_9442_), .Y(_9468_) );
	OAI21X1 OAI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_9126_), .B(_9127_), .C(_9325__bF_buf4), .Y(_9469_) );
	NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf0), .B(_9177_), .Y(_9470_) );
	OAI21X1 OAI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_9025_), .B(_9042_), .C(_9166_), .Y(_9471_) );
	AOI22X1 AOI22X1_213 ( .gnd(gnd), .vdd(vdd), .A(_9134_), .B(_9140_), .C(_9184_), .D(_9471_), .Y(_9472_) );
	OAI21X1 OAI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_9470_), .B(_9472_), .C(_9129_), .Y(_9473_) );
	INVX1 INVX1_1329 ( .gnd(gnd), .vdd(vdd), .A(_9129_), .Y(_9474_) );
	INVX1 INVX1_1330 ( .gnd(gnd), .vdd(vdd), .A(_9470_), .Y(_9475_) );
	INVX1 INVX1_1331 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .Y(_9477_) );
	NAND3X1 NAND3X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_9474_), .B(_9475_), .C(_9477_), .Y(_9478_) );
	NAND2X1 NAND2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_9473_), .B(_9478_), .Y(_9479_) );
	NAND2X1 NAND2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf3), .B(_9479_), .Y(_9480_) );
	NAND3X1 NAND3X1_2030 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf5), .B(_9469_), .C(_9480_), .Y(_9481_) );
	NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .B(divider_divuResult_2_bF_buf2), .Y(_9482_) );
	AOI21X1 AOI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_9473_), .B(_9478_), .C(_9325__bF_buf3), .Y(_9483_) );
	OAI21X1 OAI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_9483_), .C(_10678__bF_buf1), .Y(_9484_) );
	NAND2X1 NAND2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_9184_), .B(_9471_), .Y(_9485_) );
	NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(_9141_), .B(_9485_), .Y(_9486_) );
	OAI21X1 OAI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .B(_9486_), .C(divider_divuResult_2_bF_buf1), .Y(_9488_) );
	NAND2X1 NAND2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_9325__bF_buf2), .Y(_9489_) );
	NAND3X1 NAND3X1_2031 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf4), .B(_9489_), .C(_9488_), .Y(_9490_) );
	NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_9472_), .B(_9486_), .Y(_9491_) );
	NAND2X1 NAND2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_9491_), .B(divider_divuResult_2_bF_buf0), .Y(_9492_) );
	NAND3X1 NAND3X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_9132_), .B(_9133_), .C(_9325__bF_buf1), .Y(_9493_) );
	NAND3X1 NAND3X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf1), .B(_9492_), .C(_9493_), .Y(_9494_) );
	AOI22X1 AOI22X1_214 ( .gnd(gnd), .vdd(vdd), .A(_9490_), .B(_9494_), .C(_9481_), .D(_9484_), .Y(_9495_) );
	NAND2X1 NAND2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_9148_), .B(_9152_), .Y(_9496_) );
	XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9496_), .Y(_9497_) );
	OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf0), .B(_9497_), .Y(_9499_) );
	NAND3X1 NAND3X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_9150_), .B(_9151_), .C(_9325__bF_buf6), .Y(_9500_) );
	NAND3X1 NAND3X1_2035 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf2), .B(_9500_), .C(_9499_), .Y(_9501_) );
	NAND2X1 NAND2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .B(_9325__bF_buf5), .Y(_9502_) );
	NAND2X1 NAND2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(divider_divuResult_2_bF_buf7), .Y(_9503_) );
	NAND3X1 NAND3X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf1), .B(_9503_), .C(_9502_), .Y(_9504_) );
	OAI21X1 OAI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_8628_), .B(divider_divuResult_3_bF_buf7), .C(_9164_), .Y(_9505_) );
	NAND2X1 NAND2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_9505_), .B(_9325__bF_buf4), .Y(_9506_) );
	NAND2X1 NAND2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(_9165_), .Y(_9507_) );
	AOI21X1 AOI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_9299_), .B(_9496_), .C(_9181_), .Y(_9508_) );
	XNOR2X1 XNOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_9508_), .B(_9507_), .Y(_9510_) );
	NAND2X1 NAND2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_9510_), .B(divider_divuResult_2_bF_buf6), .Y(_9511_) );
	NAND2X1 NAND2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_9511_), .B(_9506_), .Y(_9512_) );
	NAND2X1 NAND2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf6), .B(_9512_), .Y(_9513_) );
	NAND3X1 NAND3X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf1), .B(_9511_), .C(_9506_), .Y(_9514_) );
	AOI22X1 AOI22X1_215 ( .gnd(gnd), .vdd(vdd), .A(_9501_), .B(_9504_), .C(_9514_), .D(_9513_), .Y(_9515_) );
	AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_9515_), .B(_9495_), .Y(_9516_) );
	NAND2X1 NAND2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_9516_), .B(_9468_), .Y(_9517_) );
	NOR3X1 NOR3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf0), .B(_9482_), .C(_9483_), .Y(_9518_) );
	AOI21X1 AOI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_9469_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf4), .Y(_9519_) );
	NAND2X1 NAND2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_9490_), .B(_9494_), .Y(_9521_) );
	OAI21X1 OAI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_9519_), .B(_9518_), .C(_9521_), .Y(_9522_) );
	NOR3X1 NOR3X1_95 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf3), .B(_9482_), .C(_9483_), .Y(_9523_) );
	OAI21X1 OAI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_9483_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf2), .Y(_9524_) );
	OAI21X1 OAI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf3), .B(_9491_), .C(_9489_), .Y(_9525_) );
	NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf3), .B(_9525_), .Y(_9526_) );
	OAI21X1 OAI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_9523_), .B(_9526_), .C(_9524_), .Y(_9527_) );
	AOI21X1 AOI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_9502_), .B(_9503_), .C(divider_absoluteValue_B_flipSign_result_7_bF_buf1), .Y(_9528_) );
	AOI21X1 AOI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_9506_), .B(_9511_), .C(divider_absoluteValue_B_flipSign_result_8_bF_buf5), .Y(_9529_) );
	NAND3X1 NAND3X1_2038 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf4), .B(_9511_), .C(_9506_), .Y(_9530_) );
	OAI21X1 OAI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_9528_), .B(_9529_), .C(_9530_), .Y(_9532_) );
	OAI21X1 OAI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_9532_), .B(_9522_), .C(_9527_), .Y(_9533_) );
	NAND2X1 NAND2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_9428_), .B(_9434_), .Y(_9534_) );
	NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf1), .B(_9440_), .Y(_9535_) );
	AOI21X1 AOI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_9438_), .B(_9437_), .C(divider_absoluteValue_B_flipSign_result_13_bF_buf1), .Y(_9536_) );
	OAI21X1 OAI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_9536_), .B(_9535_), .C(_9534_), .Y(_9537_) );
	OAI21X1 OAI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf2), .B(_9453_), .C(_9451_), .Y(_9538_) );
	NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf2), .B(_9538_), .Y(_9539_) );
	OAI21X1 OAI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_9456_), .B(_9455_), .C(divider_absoluteValue_B_flipSign_result_12_bF_buf1), .Y(_9540_) );
	AOI21X1 AOI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_9463_), .B(_9464_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf4), .Y(_9541_) );
	AOI21X1 AOI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_9541_), .C(_9539_), .Y(_9543_) );
	OAI21X1 OAI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_9313_), .B(divider_divuResult_2_bF_buf5), .C(_9427_), .Y(_9544_) );
	NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf5), .B(_9544_), .Y(_9545_) );
	NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf0), .B(_9440_), .Y(_9546_) );
	AOI21X1 AOI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_9534_), .B(_9546_), .C(_9545_), .Y(_9547_) );
	OAI21X1 OAI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_9543_), .B(_9537_), .C(_9547_), .Y(_9548_) );
	AOI21X1 AOI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .B(_9468_), .C(_9548_), .Y(_9549_) );
	OAI21X1 OAI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_9412_), .B(_9517_), .C(_9549_), .Y(_9550_) );
	OAI21X1 OAI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(divider_divuResult_2_bF_buf4), .C(_2229__bF_buf4), .Y(_9551_) );
	NAND2X1 NAND2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_30_), .B(_9551_), .Y(_9552_) );
	INVX1 INVX1_1332 ( .gnd(gnd), .vdd(vdd), .A(_9551_), .Y(_9554_) );
	NAND2X1 NAND2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_9554_), .Y(_9555_) );
	NAND2X1 NAND2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_9171_), .B(_9415_), .Y(_9556_) );
	AOI21X1 AOI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_9290_), .B(_9298_), .C(_9556_), .Y(_9557_) );
	OAI21X1 OAI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9557_), .C(_9227_), .Y(_9558_) );
	AOI21X1 AOI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_9558_), .B(_9279_), .C(_8831_), .Y(_9559_) );
	OAI21X1 OAI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .B(_9559_), .C(_8742_), .Y(_9560_) );
	AOI22X1 AOI22X1_216 ( .gnd(gnd), .vdd(vdd), .A(_8710_), .B(_8716_), .C(_9254_), .D(_9560_), .Y(_9561_) );
	NAND2X1 NAND2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_8716_), .B(_8710_), .Y(_9562_) );
	INVX1 INVX1_1333 ( .gnd(gnd), .vdd(vdd), .A(_9226_), .Y(_9563_) );
	NAND3X1 NAND3X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_8868_), .B(_8895_), .C(_9563_), .Y(_9565_) );
	AOI21X1 AOI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_9170_), .B(_9200_), .C(_9565_), .Y(_9566_) );
	OAI21X1 OAI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_8969_), .B(_9566_), .C(_9262_), .Y(_9567_) );
	AOI21X1 AOI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_9567_), .B(_8803_), .C(_8822_), .Y(_9568_) );
	NOR3X1 NOR3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .B(_8808_), .C(_9568_), .Y(_9569_) );
	OAI21X1 OAI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_9569_), .B(_9561_), .C(divider_divuResult_2_bF_buf3), .Y(_9570_) );
	OAI21X1 OAI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_8707_), .B(divider_divuResult_3_bF_buf6), .C(_8714_), .Y(_9571_) );
	OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf2), .B(_9571_), .Y(_9572_) );
	NAND3X1 NAND3X1_2040 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .B(_9572_), .C(_9570_), .Y(_9573_) );
	OAI21X1 OAI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_8808_), .B(_9568_), .C(_9562_), .Y(_9574_) );
	INVX1 INVX1_1334 ( .gnd(gnd), .vdd(vdd), .A(_9562_), .Y(_9576_) );
	NAND3X1 NAND3X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_9576_), .B(_9254_), .C(_9560_), .Y(_9577_) );
	NAND3X1 NAND3X1_2042 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf1), .B(_9574_), .C(_9577_), .Y(_9578_) );
	NAND2X1 NAND2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_9571_), .B(_9325__bF_buf1), .Y(_9579_) );
	NAND3X1 NAND3X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_9579_), .C(_9578_), .Y(_9580_) );
	AOI22X1 AOI22X1_217 ( .gnd(gnd), .vdd(vdd), .A(_9552_), .B(_9555_), .C(_9580_), .D(_9573_), .Y(_9581_) );
	OAI21X1 OAI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_8729_), .B(_8732_), .C(_9325__bF_buf0), .Y(_9582_) );
	NAND2X1 NAND2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_8728_), .B(_8733_), .Y(_9583_) );
	OAI21X1 OAI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_9251_), .B(_9559_), .C(_8821_), .Y(_9584_) );
	NAND3X1 NAND3X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_9583_), .B(_8807_), .C(_9584_), .Y(_9585_) );
	INVX1 INVX1_1335 ( .gnd(gnd), .vdd(vdd), .A(_9583_), .Y(_9587_) );
	AOI21X1 AOI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_9567_), .B(_8803_), .C(_8741_), .Y(_9588_) );
	OAI21X1 OAI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_9253_), .B(_9588_), .C(_9587_), .Y(_9589_) );
	NAND3X1 NAND3X1_2045 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf0), .B(_9589_), .C(_9585_), .Y(_9590_) );
	NAND3X1 NAND3X1_2046 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .B(_9582_), .C(_9590_), .Y(_9591_) );
	OAI21X1 OAI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_9253_), .B(_9588_), .C(_9583_), .Y(_9592_) );
	NAND3X1 NAND3X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_9587_), .B(_8807_), .C(_9584_), .Y(_9593_) );
	NAND3X1 NAND3X1_2048 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf7), .B(_9592_), .C(_9593_), .Y(_9594_) );
	NAND2X1 NAND2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_8718_), .B(_8727_), .Y(_9595_) );
	OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf6), .B(_9595_), .Y(_9596_) );
	NAND3X1 NAND3X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_9596_), .C(_9594_), .Y(_9598_) );
	OAI21X1 OAI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_9565_), .B(_9321_), .C(_9279_), .Y(_9599_) );
	AOI21X1 AOI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_9599_), .B(_9262_), .C(_9251_), .Y(_9600_) );
	AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(_8741_), .Y(_9601_) );
	OAI21X1 OAI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_9600_), .C(divider_divuResult_2_bF_buf5), .Y(_9602_) );
	NAND2X1 NAND2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_9325__bF_buf6), .Y(_9603_) );
	OAI21X1 OAI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_9601_), .B(_9602_), .C(_9603_), .Y(_9604_) );
	NAND2X1 NAND2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_9604_), .Y(_9605_) );
	NAND2X1 NAND2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_9600_), .Y(_9606_) );
	NAND3X1 NAND3X1_2050 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf4), .B(_9606_), .C(_9584_), .Y(_9607_) );
	NAND3X1 NAND3X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_9603_), .C(_9607_), .Y(_9609_) );
	AOI22X1 AOI22X1_218 ( .gnd(gnd), .vdd(vdd), .A(_9605_), .B(_9609_), .C(_9591_), .D(_9598_), .Y(_9610_) );
	NAND2X1 NAND2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_9610_), .B(_9581_), .Y(_9611_) );
	OAI21X1 OAI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_8756_), .B(divider_divuResult_3_bF_buf5), .C(_8754_), .Y(_9612_) );
	NAND2X1 NAND2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_9612_), .B(_9325__bF_buf5), .Y(_9613_) );
	NAND2X1 NAND2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_8755_), .B(_8761_), .Y(_9614_) );
	AOI21X1 AOI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_9558_), .B(_9279_), .C(_9261_), .Y(_9615_) );
	OAI21X1 OAI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_8798_), .B(_9615_), .C(_9243_), .Y(_9616_) );
	NAND3X1 NAND3X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_9614_), .B(_8801_), .C(_9616_), .Y(_9617_) );
	INVX1 INVX1_1336 ( .gnd(gnd), .vdd(vdd), .A(_9614_), .Y(_9618_) );
	OAI21X1 OAI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_8969_), .B(_9566_), .C(_8830_), .Y(_9620_) );
	AOI22X1 AOI22X1_219 ( .gnd(gnd), .vdd(vdd), .A(_8768_), .B(_8774_), .C(_9247_), .D(_9620_), .Y(_9621_) );
	OAI21X1 OAI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_9249_), .B(_9621_), .C(_9618_), .Y(_9622_) );
	NAND3X1 NAND3X1_2053 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf3), .B(_9622_), .C(_9617_), .Y(_9623_) );
	NAND3X1 NAND3X1_2054 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf2), .B(_9613_), .C(_9623_), .Y(_9624_) );
	OAI21X1 OAI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_9249_), .B(_9621_), .C(_9614_), .Y(_9625_) );
	NAND3X1 NAND3X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_9618_), .B(_8801_), .C(_9616_), .Y(_9626_) );
	NAND3X1 NAND3X1_2056 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf2), .B(_9625_), .C(_9626_), .Y(_9627_) );
	INVX1 INVX1_1337 ( .gnd(gnd), .vdd(vdd), .A(_9612_), .Y(_9628_) );
	NAND2X1 NAND2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_9628_), .B(_9325__bF_buf4), .Y(_9629_) );
	NAND3X1 NAND3X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_9629_), .C(_9627_), .Y(_9631_) );
	INVX1 INVX1_1338 ( .gnd(gnd), .vdd(vdd), .A(_9243_), .Y(_9632_) );
	AOI21X1 AOI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_9599_), .B(_8830_), .C(_8798_), .Y(_9633_) );
	AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_9633_), .B(_9632_), .Y(_9634_) );
	OAI21X1 OAI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_9632_), .B(_9633_), .C(divider_divuResult_2_bF_buf1), .Y(_9635_) );
	NAND3X1 NAND3X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_8766_), .B(_8767_), .C(_9325__bF_buf3), .Y(_9636_) );
	OAI21X1 OAI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_9634_), .B(_9635_), .C(_9636_), .Y(_9637_) );
	NAND2X1 NAND2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_9637_), .Y(_9638_) );
	NAND2X1 NAND2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_9632_), .B(_9633_), .Y(_9639_) );
	NAND3X1 NAND3X1_2059 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf0), .B(_9639_), .C(_9616_), .Y(_9640_) );
	NAND3X1 NAND3X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_9636_), .C(_9640_), .Y(_9642_) );
	AOI22X1 AOI22X1_220 ( .gnd(gnd), .vdd(vdd), .A(_9638_), .B(_9642_), .C(_9624_), .D(_9631_), .Y(_9643_) );
	OAI21X1 OAI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_8969_), .B(_9566_), .C(_9260_), .Y(_9644_) );
	OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_9599_), .B(_9260_), .Y(_9645_) );
	NAND3X1 NAND3X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_9644_), .B(_9645_), .C(divider_divuResult_2_bF_buf7), .Y(_9646_) );
	OAI21X1 OAI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_8796_), .B(divider_divuResult_2_bF_buf6), .C(_9646_), .Y(_9647_) );
	NAND2X1 NAND2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf2), .B(_9647_), .Y(_9648_) );
	OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf5), .B(_8796_), .Y(_9649_) );
	NAND3X1 NAND3X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf0), .B(_9646_), .C(_9649_), .Y(_9650_) );
	OAI21X1 OAI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_8777_), .B(_8789_), .C(_9325__bF_buf2), .Y(_9651_) );
	NAND2X1 NAND2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_8824_), .Y(_9653_) );
	NAND3X1 NAND3X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_8826_), .B(_9653_), .C(_9644_), .Y(_9654_) );
	INVX1 INVX1_1339 ( .gnd(gnd), .vdd(vdd), .A(_8826_), .Y(_9655_) );
	INVX1 INVX1_1340 ( .gnd(gnd), .vdd(vdd), .A(_9653_), .Y(_9656_) );
	AOI21X1 AOI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_9558_), .B(_9279_), .C(_8829_), .Y(_9657_) );
	OAI21X1 OAI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_9655_), .B(_9657_), .C(_9656_), .Y(_9658_) );
	NAND3X1 NAND3X1_2064 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf4), .B(_9654_), .C(_9658_), .Y(_9659_) );
	NAND3X1 NAND3X1_2065 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf1), .B(_9651_), .C(_9659_), .Y(_9660_) );
	INVX1 INVX1_1341 ( .gnd(gnd), .vdd(vdd), .A(_9651_), .Y(_9661_) );
	OAI21X1 OAI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_9655_), .B(_9657_), .C(_9653_), .Y(_9662_) );
	NAND3X1 NAND3X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_8826_), .B(_9656_), .C(_9644_), .Y(_9664_) );
	AOI21X1 AOI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_9662_), .B(_9664_), .C(_9325__bF_buf1), .Y(_9665_) );
	OAI21X1 OAI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_9661_), .B(_9665_), .C(_2042__bF_buf2), .Y(_9666_) );
	AOI22X1 AOI22X1_221 ( .gnd(gnd), .vdd(vdd), .A(_9648_), .B(_9650_), .C(_9660_), .D(_9666_), .Y(_9667_) );
	NAND2X1 NAND2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_9667_), .B(_9643_), .Y(_9668_) );
	NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_9668_), .B(_9611_), .Y(_9669_) );
	OAI21X1 OAI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_8849_), .B(divider_divuResult_3_bF_buf4), .C(_8847_), .Y(_9670_) );
	NAND2X1 NAND2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_9670_), .B(_9325__bF_buf0), .Y(_9671_) );
	NAND2X1 NAND2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_8855_), .Y(_9672_) );
	OAI21X1 OAI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9557_), .C(_9563_), .Y(_9673_) );
	AOI21X1 AOI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_9673_), .B(_8956_), .C(_9208_), .Y(_9675_) );
	OAI21X1 OAI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(_9675_), .C(_9204_), .Y(_9676_) );
	NAND3X1 NAND3X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_9672_), .B(_8966_), .C(_9676_), .Y(_9677_) );
	INVX1 INVX1_1342 ( .gnd(gnd), .vdd(vdd), .A(_9672_), .Y(_9678_) );
	AOI21X1 AOI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_9170_), .B(_9200_), .C(_9226_), .Y(_9679_) );
	OAI21X1 OAI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_9271_), .B(_9679_), .C(_8895_), .Y(_9680_) );
	AOI22X1 AOI22X1_222 ( .gnd(gnd), .vdd(vdd), .A(_8863_), .B(_8867_), .C(_9274_), .D(_9680_), .Y(_9681_) );
	OAI21X1 OAI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_8965_), .B(_9681_), .C(_9678_), .Y(_9682_) );
	NAND3X1 NAND3X1_2068 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf3), .B(_9682_), .C(_9677_), .Y(_9683_) );
	NAND3X1 NAND3X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf2), .B(_9671_), .C(_9683_), .Y(_9684_) );
	INVX1 INVX1_1343 ( .gnd(gnd), .vdd(vdd), .A(_9670_), .Y(_9686_) );
	NAND2X1 NAND2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_9686_), .B(_9325__bF_buf6), .Y(_9687_) );
	OAI21X1 OAI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_8965_), .B(_9681_), .C(_9672_), .Y(_9688_) );
	NAND3X1 NAND3X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_9678_), .B(_8966_), .C(_9676_), .Y(_9689_) );
	NAND3X1 NAND3X1_2071 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf2), .B(_9688_), .C(_9689_), .Y(_9690_) );
	NAND3X1 NAND3X1_2072 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf0), .B(_9687_), .C(_9690_), .Y(_9691_) );
	INVX1 INVX1_1344 ( .gnd(gnd), .vdd(vdd), .A(_9204_), .Y(_9692_) );
	INVX1 INVX1_1345 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .Y(_9693_) );
	OAI21X1 OAI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf4), .B(_9693_), .C(_8957_), .Y(_9694_) );
	OAI21X1 OAI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_9226_), .B(_9321_), .C(_8956_), .Y(_9695_) );
	AOI22X1 AOI22X1_223 ( .gnd(gnd), .vdd(vdd), .A(_9206_), .B(_9694_), .C(_8895_), .D(_9695_), .Y(_9697_) );
	AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_9697_), .B(_9692_), .Y(_9698_) );
	OAI21X1 OAI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_9692_), .B(_9697_), .C(divider_divuResult_2_bF_buf1), .Y(_9699_) );
	NAND3X1 NAND3X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_8859_), .B(_8862_), .C(_9325__bF_buf5), .Y(_9700_) );
	OAI21X1 OAI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_9698_), .B(_9699_), .C(_9700_), .Y(_9701_) );
	NAND2X1 NAND2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf0), .B(_9701_), .Y(_9702_) );
	NAND2X1 NAND2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_9692_), .B(_9697_), .Y(_9703_) );
	NAND3X1 NAND3X1_2074 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf0), .B(_9703_), .C(_9676_), .Y(_9704_) );
	NAND3X1 NAND3X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf0), .B(_9700_), .C(_9704_), .Y(_9705_) );
	NAND2X1 NAND2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_9705_), .B(_9702_), .Y(_9706_) );
	NAND3X1 NAND3X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_9684_), .B(_9691_), .C(_9706_), .Y(_9708_) );
	OAI21X1 OAI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(divider_divuResult_3_bF_buf3), .C(_8877_), .Y(_9709_) );
	NAND2X1 NAND2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_9709_), .B(_9325__bF_buf4), .Y(_9710_) );
	NAND2X1 NAND2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_8885_), .B(_8878_), .Y(_9711_) );
	OAI21X1 OAI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_9271_), .B(_9679_), .C(_9207_), .Y(_9712_) );
	NAND3X1 NAND3X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_9711_), .B(_8961_), .C(_9712_), .Y(_9713_) );
	INVX1 INVX1_1346 ( .gnd(gnd), .vdd(vdd), .A(_9207_), .Y(_9714_) );
	AOI21X1 AOI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .B(_9563_), .C(_9271_), .Y(_9715_) );
	OAI21X1 OAI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_9714_), .B(_9715_), .C(_8961_), .Y(_9716_) );
	OAI21X1 OAI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_9272_), .B(_8958_), .C(_9716_), .Y(_9717_) );
	NAND3X1 NAND3X1_2078 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf7), .B(_9713_), .C(_9717_), .Y(_9719_) );
	NAND3X1 NAND3X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf2), .B(_9710_), .C(_9719_), .Y(_9720_) );
	INVX1 INVX1_1347 ( .gnd(gnd), .vdd(vdd), .A(_9709_), .Y(_9721_) );
	NAND2X1 NAND2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_9721_), .B(_9325__bF_buf3), .Y(_9722_) );
	AOI21X1 AOI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_8878_), .B(_8885_), .C(_9716_), .Y(_9723_) );
	AOI21X1 AOI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_9712_), .B(_8961_), .C(_9711_), .Y(_9724_) );
	OAI21X1 OAI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_9724_), .B(_9723_), .C(divider_divuResult_2_bF_buf6), .Y(_9725_) );
	NAND3X1 NAND3X1_2080 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf3), .B(_9722_), .C(_9725_), .Y(_9726_) );
	NAND2X1 NAND2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_9714_), .B(_9715_), .Y(_9727_) );
	NAND2X1 NAND2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_9712_), .B(_9727_), .Y(_9728_) );
	NAND2X1 NAND2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf5), .B(_9728_), .Y(_9730_) );
	NAND2X1 NAND2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_9693_), .B(_9325__bF_buf2), .Y(_9731_) );
	NAND3X1 NAND3X1_2081 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf3), .B(_9731_), .C(_9730_), .Y(_9732_) );
	NAND3X1 NAND3X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_9712_), .B(_9727_), .C(divider_divuResult_2_bF_buf4), .Y(_9733_) );
	NAND2X1 NAND2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(_9325__bF_buf1), .Y(_9734_) );
	NAND3X1 NAND3X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf0), .B(_9734_), .C(_9733_), .Y(_9735_) );
	NAND2X1 NAND2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_9735_), .B(_9732_), .Y(_9736_) );
	NAND3X1 NAND3X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_9720_), .B(_9736_), .C(_9726_), .Y(_9737_) );
	NAND2X1 NAND2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .B(_9325__bF_buf0), .Y(_9738_) );
	NAND2X1 NAND2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .B(_9219_), .Y(_9739_) );
	NAND2X1 NAND2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_9223_), .B(_9222_), .Y(_9741_) );
	NAND2X1 NAND2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_9741_), .B(_9739_), .Y(_9742_) );
	AOI21X1 AOI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_9170_), .B(_9200_), .C(_9742_), .Y(_9743_) );
	OAI21X1 OAI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_8954_), .B(_9743_), .C(_9212_), .Y(_9744_) );
	NAND3X1 NAND3X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_9211_), .B(_8923_), .C(_9744_), .Y(_9745_) );
	INVX1 INVX1_1348 ( .gnd(gnd), .vdd(vdd), .A(_8954_), .Y(_9746_) );
	OAI21X1 OAI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9557_), .C(_9225_), .Y(_9747_) );
	AOI21X1 AOI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_9747_), .B(_9746_), .C(_8931_), .Y(_9748_) );
	OAI21X1 OAI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_9269_), .B(_9748_), .C(_8919_), .Y(_9749_) );
	NAND3X1 NAND3X1_2086 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf3), .B(_9745_), .C(_9749_), .Y(_9750_) );
	NAND3X1 NAND3X1_2087 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf3), .B(_9738_), .C(_9750_), .Y(_9752_) );
	OAI21X1 OAI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_9269_), .B(_9748_), .C(_9211_), .Y(_9753_) );
	NAND3X1 NAND3X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_8919_), .B(_8923_), .C(_9744_), .Y(_9754_) );
	NAND3X1 NAND3X1_2089 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf2), .B(_9754_), .C(_9753_), .Y(_9755_) );
	NAND2X1 NAND2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .B(_9325__bF_buf6), .Y(_9756_) );
	NAND3X1 NAND3X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf2), .B(_9756_), .C(_9755_), .Y(_9757_) );
	NAND2X1 NAND2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_9752_), .B(_9757_), .Y(_9758_) );
	NAND3X1 NAND3X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_9746_), .C(_9747_), .Y(_9759_) );
	NAND2X1 NAND2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_9744_), .B(_9759_), .Y(_9760_) );
	NAND2X1 NAND2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf1), .B(_9760_), .Y(_9761_) );
	OAI21X1 OAI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .B(divider_divuResult_3_bF_buf2), .C(_8921_), .Y(_9763_) );
	NAND2X1 NAND2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_9763_), .B(_9325__bF_buf5), .Y(_9764_) );
	NAND3X1 NAND3X1_2092 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf3), .B(_9764_), .C(_9761_), .Y(_9765_) );
	NAND3X1 NAND3X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_9744_), .B(_9759_), .C(divider_divuResult_2_bF_buf0), .Y(_9766_) );
	INVX1 INVX1_1349 ( .gnd(gnd), .vdd(vdd), .A(_9763_), .Y(_9767_) );
	NAND2X1 NAND2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_9767_), .B(_9325__bF_buf4), .Y(_9768_) );
	NAND3X1 NAND3X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf1), .B(_9768_), .C(_9766_), .Y(_9769_) );
	NAND2X1 NAND2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_9769_), .Y(_9770_) );
	INVX1 INVX1_1350 ( .gnd(gnd), .vdd(vdd), .A(_8952_), .Y(_9771_) );
	AOI21X1 AOI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_9222_), .B(_9223_), .C(_9321_), .Y(_9772_) );
	OAI21X1 OAI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_9771_), .B(_9772_), .C(_9739_), .Y(_9774_) );
	INVX1 INVX1_1351 ( .gnd(gnd), .vdd(vdd), .A(_9739_), .Y(_9775_) );
	OAI21X1 OAI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_9557_), .C(_9741_), .Y(_9776_) );
	NAND3X1 NAND3X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_8952_), .B(_9775_), .C(_9776_), .Y(_9777_) );
	NAND2X1 NAND2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_9777_), .B(_9774_), .Y(_9778_) );
	NAND2X1 NAND2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf7), .B(_9778_), .Y(_9779_) );
	OAI21X1 OAI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_9217_), .B(_9218_), .C(_9325__bF_buf3), .Y(_9780_) );
	NAND3X1 NAND3X1_2096 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf3), .B(_9780_), .C(_9779_), .Y(_9781_) );
	AOI21X1 AOI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_9774_), .B(_9777_), .C(_9325__bF_buf2), .Y(_9782_) );
	OAI21X1 OAI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_9216_), .B(divider_divuResult_3_bF_buf1), .C(_8944_), .Y(_9783_) );
	INVX1 INVX1_1352 ( .gnd(gnd), .vdd(vdd), .A(_9783_), .Y(_9785_) );
	NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_9785_), .B(divider_divuResult_2_bF_buf6), .Y(_9786_) );
	OAI21X1 OAI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_9786_), .B(_9782_), .C(_2922__bF_buf0), .Y(_9787_) );
	NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_9741_), .B(_9201_), .Y(_9788_) );
	OAI21X1 OAI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_9772_), .B(_9788_), .C(divider_divuResult_2_bF_buf5), .Y(_9789_) );
	NAND3X1 NAND3X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_8946_), .B(_8950_), .C(_9325__bF_buf1), .Y(_9790_) );
	NAND3X1 NAND3X1_2098 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf3), .B(_9789_), .C(_9790_), .Y(_9791_) );
	NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_9772_), .B(_9788_), .Y(_9792_) );
	NAND2X1 NAND2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_9792_), .B(divider_divuResult_2_bF_buf4), .Y(_9793_) );
	NAND2X1 NAND2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(_9325__bF_buf0), .Y(_9794_) );
	NAND3X1 NAND3X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf2), .B(_9793_), .C(_9794_), .Y(_9796_) );
	AOI22X1 AOI22X1_224 ( .gnd(gnd), .vdd(vdd), .A(_9791_), .B(_9796_), .C(_9781_), .D(_9787_), .Y(_9797_) );
	NAND3X1 NAND3X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_9770_), .B(_9797_), .C(_9758_), .Y(_9798_) );
	NOR3X1 NOR3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .B(_9798_), .C(_9708_), .Y(_9799_) );
	NAND3X1 NAND3X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_9799_), .B(_9669_), .C(_9550_), .Y(_9800_) );
	NAND3X1 NAND3X1_2102 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf3), .B(_9671_), .C(_9683_), .Y(_9801_) );
	NAND3X1 NAND3X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf1), .B(_9687_), .C(_9690_), .Y(_9802_) );
	AOI22X1 AOI22X1_225 ( .gnd(gnd), .vdd(vdd), .A(_9702_), .B(_9705_), .C(_9801_), .D(_9802_), .Y(_9803_) );
	INVX1 INVX1_1353 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .Y(_9804_) );
	NAND3X1 NAND3X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf1), .B(_9738_), .C(_9750_), .Y(_9805_) );
	NAND3X1 NAND3X1_2105 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf2), .B(_9756_), .C(_9755_), .Y(_9807_) );
	NAND3X1 NAND3X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_9805_), .B(_9807_), .C(_9770_), .Y(_9808_) );
	NOR3X1 NOR3X1_98 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf2), .B(_9786_), .C(_9782_), .Y(_9809_) );
	OAI21X1 OAI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_9786_), .B(_9782_), .C(divider_absoluteValue_B_flipSign_result_16_bF_buf1), .Y(_9810_) );
	AOI21X1 AOI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_9794_), .B(_9793_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf2), .Y(_9811_) );
	OAI21X1 OAI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_9811_), .B(_9809_), .C(_9810_), .Y(_9812_) );
	AOI21X1 AOI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_9755_), .B(_9756_), .C(divider_absoluteValue_B_flipSign_result_18_bF_buf1), .Y(_9813_) );
	OAI21X1 OAI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_9767_), .B(divider_divuResult_2_bF_buf3), .C(_9761_), .Y(_9814_) );
	NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf2), .B(_9814_), .Y(_9815_) );
	AOI21X1 AOI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_9815_), .B(_9807_), .C(_9813_), .Y(_9816_) );
	OAI21X1 OAI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_9812_), .B(_9808_), .C(_9816_), .Y(_9818_) );
	NAND3X1 NAND3X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_9803_), .B(_9804_), .C(_9818_), .Y(_9819_) );
	OAI21X1 OAI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf6), .B(_9728_), .C(_9734_), .Y(_9820_) );
	NAND2X1 NAND2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf4), .B(_9820_), .Y(_9821_) );
	NAND2X1 NAND2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_9821_), .B(_9720_), .Y(_9822_) );
	AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_9822_), .B(_9726_), .Y(_9823_) );
	NAND2X1 NAND2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_9803_), .B(_9823_), .Y(_9824_) );
	AOI21X1 AOI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_9690_), .B(_9687_), .C(divider_absoluteValue_B_flipSign_result_22_bF_buf2), .Y(_9825_) );
	NAND2X1 NAND2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf3), .B(_9701_), .Y(_9826_) );
	INVX1 INVX1_1354 ( .gnd(gnd), .vdd(vdd), .A(_9826_), .Y(_9827_) );
	AOI21X1 AOI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_9827_), .B(_9691_), .C(_9825_), .Y(_9829_) );
	NAND3X1 NAND3X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_9824_), .B(_9829_), .C(_9819_), .Y(_9830_) );
	NAND2X1 NAND2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf3), .B(_9647_), .Y(_9831_) );
	NAND3X1 NAND3X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf1), .B(_9651_), .C(_9659_), .Y(_9832_) );
	AOI21X1 AOI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_9659_), .B(_9651_), .C(_2042__bF_buf0), .Y(_9833_) );
	AOI21X1 AOI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_9831_), .B(_9832_), .C(_9833_), .Y(_9834_) );
	NAND3X1 NAND3X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_9613_), .C(_9623_), .Y(_9835_) );
	AOI21X1 AOI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_9623_), .B(_9613_), .C(_6845_), .Y(_9836_) );
	NAND2X1 NAND2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_9637_), .Y(_9837_) );
	OAI21X1 OAI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_9837_), .B(_9836_), .C(_9835_), .Y(_9838_) );
	AOI21X1 AOI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_9643_), .B(_9834_), .C(_9838_), .Y(_9840_) );
	NAND3X1 NAND3X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_9582_), .C(_9590_), .Y(_9841_) );
	AOI21X1 AOI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_9590_), .B(_9582_), .C(_2009_), .Y(_9842_) );
	NAND2X1 NAND2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_9604_), .Y(_9843_) );
	OAI21X1 OAI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .B(_9842_), .C(_9841_), .Y(_9844_) );
	NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_30_), .B(_9554_), .Y(_9845_) );
	INVX1 INVX1_1355 ( .gnd(gnd), .vdd(vdd), .A(_9845_), .Y(_9846_) );
	NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_9551_), .Y(_9847_) );
	NAND3X1 NAND3X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_9572_), .C(_9570_), .Y(_9848_) );
	OAI21X1 OAI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_9847_), .B(_9848_), .C(_9846_), .Y(_9849_) );
	AOI21X1 AOI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_9581_), .B(_9844_), .C(_9849_), .Y(_9851_) );
	OAI21X1 OAI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_9611_), .B(_9840_), .C(_9851_), .Y(_9852_) );
	AOI21X1 AOI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_9669_), .B(_9830_), .C(_9852_), .Y(_9853_) );
	AOI21X1 AOI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_9853_), .B(_9800_), .C(divider_absoluteValue_B_flipSign_result_31_), .Y(divider_divuResult_1_) );
	OAI21X1 OAI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_9686_), .B(divider_divuResult_2_bF_buf2), .C(_9683_), .Y(_9854_) );
	AOI21X1 AOI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_9328_), .B(_9332_), .C(_9239_), .Y(_9855_) );
	INVX1 INVX1_1356 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_2_), .Y(_9856_) );
	NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf3), .B(_9856_), .Y(_9857_) );
	NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_9857_), .Y(_9858_) );
	NAND2X1 NAND2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_9858_), .B(divider_divuResult_2_bF_buf1), .Y(_9859_) );
	NAND2X1 NAND2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_9856_), .B(_9325__bF_buf5), .Y(_9861_) );
	NAND3X1 NAND3X1_2113 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf0), .B(_9859_), .C(_9861_), .Y(_9862_) );
	NAND3X1 NAND3X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf4), .B(_9331_), .C(_9330_), .Y(_9863_) );
	NAND2X1 NAND2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_9862_), .B(_9863_), .Y(_9864_) );
	NAND3X1 NAND3X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_8586_), .B(_8660_), .C(_9325__bF_buf4), .Y(_9865_) );
	NAND3X1 NAND3X1_2116 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf2), .B(_9237_), .C(_9865_), .Y(_9866_) );
	OAI21X1 OAI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9326_), .C(_2547__bF_buf4), .Y(_9867_) );
	NAND2X1 NAND2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_9866_), .B(_9867_), .Y(_9868_) );
	NAND3X1 NAND3X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .B(_9864_), .C(_9868_), .Y(_9869_) );
	NAND2X1 NAND2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_9363_), .B(_9393_), .Y(_9870_) );
	AOI21X1 AOI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_9869_), .B(_9855_), .C(_9870_), .Y(_9872_) );
	NAND2X1 NAND2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_9442_), .B(_9467_), .Y(_9873_) );
	NAND2X1 NAND2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_9515_), .Y(_9874_) );
	NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_9874_), .B(_9873_), .Y(_9875_) );
	OAI21X1 OAI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9872_), .C(_9875_), .Y(_9876_) );
	NAND2X1 NAND2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_9552_), .B(_9555_), .Y(_9877_) );
	NAND3X1 NAND3X1_2118 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .B(_9579_), .C(_9578_), .Y(_9878_) );
	NAND3X1 NAND3X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_9877_), .B(_9878_), .C(_9848_), .Y(_9879_) );
	NAND3X1 NAND3X1_2120 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .B(_9596_), .C(_9594_), .Y(_9880_) );
	NAND2X1 NAND2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_9609_), .B(_9605_), .Y(_9881_) );
	NAND3X1 NAND3X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_9841_), .B(_9880_), .C(_9881_), .Y(_9883_) );
	NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_9883_), .B(_9879_), .Y(_9884_) );
	AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_9643_), .B(_9667_), .Y(_9885_) );
	NAND3X1 NAND3X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_9885_), .B(_9884_), .C(_9799_), .Y(_9886_) );
	AOI21X1 AOI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_9876_), .B(_9549_), .C(_9886_), .Y(_9887_) );
	NAND2X1 NAND2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_9885_), .B(_9884_), .Y(_9888_) );
	NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .B(_9708_), .Y(_9889_) );
	OAI21X1 OAI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_9721_), .B(divider_divuResult_2_bF_buf0), .C(_9719_), .Y(_9890_) );
	INVX1 INVX1_1357 ( .gnd(gnd), .vdd(vdd), .A(_9890_), .Y(_9891_) );
	OAI21X1 OAI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf1), .B(_9891_), .C(_9822_), .Y(_9892_) );
	OAI21X1 OAI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_9892_), .B(_9708_), .C(_9829_), .Y(_9894_) );
	AOI21X1 AOI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_9889_), .B(_9818_), .C(_9894_), .Y(_9895_) );
	NAND3X1 NAND3X1_2123 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf1), .B(_9629_), .C(_9627_), .Y(_9896_) );
	NAND2X1 NAND2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_9642_), .B(_9638_), .Y(_9897_) );
	NAND3X1 NAND3X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_9835_), .B(_9896_), .C(_9897_), .Y(_9898_) );
	INVX1 INVX1_1358 ( .gnd(gnd), .vdd(vdd), .A(_9834_), .Y(_9899_) );
	AOI21X1 AOI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_9627_), .B(_9629_), .C(divider_absoluteValue_B_flipSign_result_26_bF_buf0), .Y(_9900_) );
	INVX1 INVX1_1359 ( .gnd(gnd), .vdd(vdd), .A(_9837_), .Y(_9901_) );
	AOI21X1 AOI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_9901_), .B(_9896_), .C(_9900_), .Y(_9902_) );
	OAI21X1 OAI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_9899_), .B(_9898_), .C(_9902_), .Y(_9903_) );
	AOI21X1 AOI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_9594_), .B(_9596_), .C(divider_absoluteValue_B_flipSign_result_28_), .Y(_9905_) );
	INVX1 INVX1_1360 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .Y(_9906_) );
	AOI21X1 AOI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_9906_), .B(_9880_), .C(_9905_), .Y(_9907_) );
	AOI21X1 AOI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_9578_), .B(_9579_), .C(divider_absoluteValue_B_flipSign_result_29_), .Y(_9908_) );
	AOI21X1 AOI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_9908_), .B(_9877_), .C(_9845_), .Y(_9909_) );
	OAI21X1 OAI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_9907_), .B(_9879_), .C(_9909_), .Y(_9910_) );
	AOI21X1 AOI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_9884_), .B(_9903_), .C(_9910_), .Y(_9911_) );
	OAI21X1 OAI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_9888_), .B(_9895_), .C(_9911_), .Y(_9912_) );
	OAI21X1 OAI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_9887_), .B(_9912_), .C(_1560__bF_buf2), .Y(_9913_) );
	NAND2X1 NAND2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_9854_), .B(_9913__bF_buf5), .Y(_9914_) );
	NAND2X1 NAND2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_9801_), .B(_9802_), .Y(_9916_) );
	INVX1 INVX1_1361 ( .gnd(gnd), .vdd(vdd), .A(_9798_), .Y(_9917_) );
	AOI21X1 AOI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_9550_), .B(_9917_), .C(_9818_), .Y(_9918_) );
	OAI21X1 OAI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .B(_9918_), .C(_9892_), .Y(_9919_) );
	NAND2X1 NAND2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .B(_9919_), .Y(_9920_) );
	NAND3X1 NAND3X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_9916_), .B(_9826_), .C(_9920_), .Y(_9921_) );
	INVX1 INVX1_1362 ( .gnd(gnd), .vdd(vdd), .A(_9916_), .Y(_9922_) );
	AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_9919_), .B(_9706_), .Y(_9923_) );
	OAI21X1 OAI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_9827_), .B(_9923_), .C(_9922_), .Y(_9924_) );
	NAND3X1 NAND3X1_2126 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf6), .B(_9921_), .C(_9924_), .Y(_9925_) );
	NAND3X1 NAND3X1_2127 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf1), .B(_9914_), .C(_9925_), .Y(_9927_) );
	INVX1 INVX1_1363 ( .gnd(gnd), .vdd(vdd), .A(_9854_), .Y(_9928_) );
	NAND2X1 NAND2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_9928_), .B(_9913__bF_buf4), .Y(_9929_) );
	OAI21X1 OAI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_9827_), .B(_9923_), .C(_9916_), .Y(_9930_) );
	NAND3X1 NAND3X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_9922_), .B(_9826_), .C(_9920_), .Y(_9931_) );
	NAND3X1 NAND3X1_2129 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf5), .B(_9931_), .C(_9930_), .Y(_9932_) );
	NAND3X1 NAND3X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf2), .B(_9929_), .C(_9932_), .Y(_9933_) );
	NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .B(_9919_), .Y(_9934_) );
	NAND2X1 NAND2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf4), .B(_9920_), .Y(_9935_) );
	NAND2X1 NAND2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_9701_), .B(_9913__bF_buf3), .Y(_9936_) );
	OAI21X1 OAI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_9935_), .C(_9936_), .Y(_9938_) );
	NAND2X1 NAND2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_22_bF_buf1), .B(_9938_), .Y(_9939_) );
	INVX1 INVX1_1364 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .Y(_9940_) );
	NAND3X1 NAND3X1_2131 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf3), .B(_9920_), .C(_9940_), .Y(_9941_) );
	NAND3X1 NAND3X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf0), .B(_9936_), .C(_9941_), .Y(_9942_) );
	AOI22X1 AOI22X1_226 ( .gnd(gnd), .vdd(vdd), .A(_9939_), .B(_9942_), .C(_9927_), .D(_9933_), .Y(_9943_) );
	NAND2X1 NAND2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_9890_), .B(_9913__bF_buf2), .Y(_9944_) );
	NAND3X1 NAND3X1_2133 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf2), .B(_9710_), .C(_9719_), .Y(_9945_) );
	NAND2X1 NAND2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf0), .B(_9890_), .Y(_9946_) );
	NAND2X1 NAND2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_9945_), .B(_9946_), .Y(_9947_) );
	INVX1 INVX1_1365 ( .gnd(gnd), .vdd(vdd), .A(_9736_), .Y(_9949_) );
	OAI21X1 OAI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_9949_), .B(_9918_), .C(_9821_), .Y(_9950_) );
	AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_9950_), .B(_9947_), .Y(_9951_) );
	NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_9947_), .B(_9950_), .Y(_9952_) );
	OAI21X1 OAI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_9952_), .B(_9951_), .C(divider_divuResult_1_bF_buf2), .Y(_9953_) );
	NAND3X1 NAND3X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf2), .B(_9944_), .C(_9953_), .Y(_9954_) );
	OAI21X1 OAI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_9891_), .B(divider_divuResult_1_bF_buf1), .C(_9953_), .Y(_9955_) );
	NAND2X1 NAND2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_21_bF_buf3), .B(_9955_), .Y(_9956_) );
	XNOR2X1 XNOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_9918_), .B(_9949_), .Y(_9957_) );
	NAND2X1 NAND2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_9820_), .B(_9913__bF_buf1), .Y(_9958_) );
	OAI21X1 OAI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_9913__bF_buf0), .B(_9957_), .C(_9958_), .Y(_9960_) );
	XNOR2X1 XNOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_9960_), .B(divider_absoluteValue_B_flipSign_result_20_bF_buf1), .Y(_9961_) );
	NAND3X1 NAND3X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_9954_), .B(_9961_), .C(_9956_), .Y(_9962_) );
	INVX1 INVX1_1366 ( .gnd(gnd), .vdd(vdd), .A(_9962_), .Y(_9963_) );
	NAND2X1 NAND2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_9963_), .Y(_9964_) );
	OAI21X1 OAI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .B(divider_divuResult_2_bF_buf7), .C(_9755_), .Y(_9965_) );
	OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf0), .B(_9965_), .Y(_9966_) );
	INVX1 INVX1_1367 ( .gnd(gnd), .vdd(vdd), .A(_9815_), .Y(_9967_) );
	INVX1 INVX1_1368 ( .gnd(gnd), .vdd(vdd), .A(_9770_), .Y(_9968_) );
	INVX1 INVX1_1369 ( .gnd(gnd), .vdd(vdd), .A(_9812_), .Y(_9969_) );
	AOI21X1 AOI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_9550_), .B(_9797_), .C(_9969_), .Y(_9970_) );
	OAI21X1 OAI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_9968_), .B(_9970_), .C(_9967_), .Y(_9971_) );
	AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_9971_), .B(_9758_), .Y(_9972_) );
	NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_9758_), .B(_9971_), .Y(_9973_) );
	OAI21X1 OAI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_9973_), .B(_9972_), .C(divider_divuResult_1_bF_buf6), .Y(_9974_) );
	NAND3X1 NAND3X1_2136 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_19_bF_buf2), .B(_9966_), .C(_9974_), .Y(_9975_) );
	NAND2X1 NAND2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_9965_), .B(_9913__bF_buf5), .Y(_9976_) );
	INVX1 INVX1_1370 ( .gnd(gnd), .vdd(vdd), .A(_9758_), .Y(_9977_) );
	NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_9977_), .B(_9971_), .Y(_9978_) );
	AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_9971_), .B(_9977_), .Y(_9979_) );
	OAI21X1 OAI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_9978_), .B(_9979_), .C(divider_divuResult_1_bF_buf5), .Y(_9982_) );
	NAND3X1 NAND3X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf3), .B(_9976_), .C(_9982_), .Y(_9983_) );
	OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_9970_), .B(_9968_), .Y(_9984_) );
	NAND2X1 NAND2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_9968_), .B(_9970_), .Y(_9985_) );
	NAND3X1 NAND3X1_2138 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf4), .B(_9985_), .C(_9984_), .Y(_9986_) );
	OAI21X1 OAI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_9814_), .B(divider_divuResult_1_bF_buf3), .C(_9986_), .Y(_9987_) );
	NAND2X1 NAND2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_3263__bF_buf0), .B(_9987_), .Y(_9988_) );
	OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf2), .B(_9814_), .Y(_9989_) );
	NAND3X1 NAND3X1_2139 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_18_bF_buf0), .B(_9986_), .C(_9989_), .Y(_9990_) );
	NAND2X1 NAND2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_9990_), .B(_9988_), .Y(_9991_) );
	AOI21X1 AOI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_9975_), .B(_9983_), .C(_9991_), .Y(_9993_) );
	OAI21X1 OAI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_9785_), .B(divider_divuResult_2_bF_buf6), .C(_9779_), .Y(_9994_) );
	NAND2X1 NAND2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_9781_), .B(_9787_), .Y(_9995_) );
	NAND2X1 NAND2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_9796_), .B(_9791_), .Y(_9996_) );
	AOI21X1 AOI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_9550_), .B(_9996_), .C(_9811_), .Y(_9997_) );
	AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_9997_), .B(_9995_), .Y(_9998_) );
	NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_9995_), .B(_9997_), .Y(_9999_) );
	OAI21X1 OAI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_9999_), .B(_9998_), .C(divider_divuResult_1_bF_buf1), .Y(_10000_) );
	OAI21X1 OAI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_9994_), .B(divider_divuResult_1_bF_buf0), .C(_10000_), .Y(_10001_) );
	NAND2X1 NAND2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_2887__bF_buf0), .B(_10001_), .Y(_10002_) );
	OAI21X1 OAI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(divider_divuResult_2_bF_buf5), .C(_9789_), .Y(_10004_) );
	NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_10004_), .B(divider_divuResult_1_bF_buf6), .Y(_10005_) );
	XNOR2X1 XNOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_9550_), .B(_9996_), .Y(_10006_) );
	NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_10006_), .B(_9913__bF_buf4), .Y(_10007_) );
	OAI21X1 OAI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_10007_), .B(_10005_), .C(_2922__bF_buf3), .Y(_10008_) );
	OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf5), .B(_9994_), .Y(_10009_) );
	NAND3X1 NAND3X1_2140 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_17_bF_buf1), .B(_10000_), .C(_10009_), .Y(_10010_) );
	NAND2X1 NAND2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_10010_), .B(_10002_), .Y(_10011_) );
	OAI21X1 OAI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_10008_), .B(_10011_), .C(_10002_), .Y(_10012_) );
	NAND3X1 NAND3X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_3789__bF_buf2), .B(_9966_), .C(_9974_), .Y(_10013_) );
	AOI21X1 AOI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_9974_), .B(_9966_), .C(_3789__bF_buf1), .Y(_10015_) );
	OAI21X1 OAI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_9988_), .B(_10015_), .C(_10013_), .Y(_10016_) );
	AOI21X1 AOI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_10012_), .B(_9993_), .C(_10016_), .Y(_10017_) );
	INVX1 INVX1_1371 ( .gnd(gnd), .vdd(vdd), .A(_9960_), .Y(_10018_) );
	OAI21X1 OAI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_20_bF_buf0), .B(_10018_), .C(_9954_), .Y(_10019_) );
	NAND2X1 NAND2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_9956_), .B(_10019_), .Y(_10020_) );
	INVX1 INVX1_1372 ( .gnd(gnd), .vdd(vdd), .A(_10020_), .Y(_10021_) );
	NAND3X1 NAND3X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_5516__bF_buf1), .B(_9914_), .C(_9925_), .Y(_10022_) );
	NAND3X1 NAND3X1_2143 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_23_bF_buf0), .B(_9929_), .C(_9932_), .Y(_10023_) );
	NAND2X1 NAND2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_4881__bF_buf3), .B(_9938_), .Y(_10024_) );
	INVX1 INVX1_1373 ( .gnd(gnd), .vdd(vdd), .A(_10024_), .Y(_10026_) );
	NAND2X1 NAND2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_10023_), .B(_10026_), .Y(_10027_) );
	NAND2X1 NAND2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_10022_), .B(_10027_), .Y(_10028_) );
	AOI21X1 AOI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_10021_), .C(_10028_), .Y(_10029_) );
	OAI21X1 OAI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_10017_), .B(_9964_), .C(_10029_), .Y(_10030_) );
	OAI21X1 OAI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_9628_), .B(divider_divuResult_2_bF_buf4), .C(_9623_), .Y(_10031_) );
	NAND2X1 NAND2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_10031_), .B(_9913__bF_buf3), .Y(_10032_) );
	NAND2X1 NAND2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_9624_), .B(_9631_), .Y(_10033_) );
	INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(_9897_), .Y(_10034_) );
	AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_9550_), .B(_9799_), .Y(_10035_) );
	OAI21X1 OAI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .B(_10035_), .C(_9667_), .Y(_10037_) );
	AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_10037_), .B(_9899_), .Y(_10038_) );
	OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_10034_), .Y(_10039_) );
	NAND3X1 NAND3X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_10033_), .B(_9837_), .C(_10039_), .Y(_10040_) );
	OAI21X1 OAI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_10034_), .B(_10038_), .C(_9837_), .Y(_10041_) );
	OAI21X1 OAI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_9900_), .B(_9836_), .C(_10041_), .Y(_10042_) );
	NAND3X1 NAND3X1_2145 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf4), .B(_10042_), .C(_10040_), .Y(_10043_) );
	NAND3X1 NAND3X1_2146 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_27_), .B(_10032_), .C(_10043_), .Y(_10044_) );
	INVX1 INVX1_1374 ( .gnd(gnd), .vdd(vdd), .A(_10031_), .Y(_10045_) );
	NAND2X1 NAND2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_10045_), .B(_9913__bF_buf2), .Y(_10046_) );
	NAND2X1 NAND2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_10033_), .B(_10041_), .Y(_10048_) );
	OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_10041_), .B(_10033_), .Y(_10049_) );
	NAND3X1 NAND3X1_2147 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf3), .B(_10048_), .C(_10049_), .Y(_10050_) );
	NAND3X1 NAND3X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_10046_), .C(_10050_), .Y(_10051_) );
	AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_10034_), .Y(_10052_) );
	OAI21X1 OAI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_10034_), .B(_10038_), .C(divider_divuResult_1_bF_buf2), .Y(_10053_) );
	NAND2X1 NAND2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_9637_), .B(_9913__bF_buf1), .Y(_10054_) );
	OAI21X1 OAI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_10052_), .B(_10053_), .C(_10054_), .Y(_10055_) );
	NAND2X1 NAND2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_26_bF_buf3), .B(_10055_), .Y(_10056_) );
	OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_10055_), .B(divider_absoluteValue_B_flipSign_result_26_bF_buf2), .Y(_10057_) );
	AOI22X1 AOI22X1_227 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_10057_), .C(_10044_), .D(_10051_), .Y(_10059_) );
	OAI21X1 OAI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_9661_), .B(_9665_), .C(_9913__bF_buf0), .Y(_10060_) );
	NAND2X1 NAND2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_9660_), .B(_9666_), .Y(_10061_) );
	INVX1 INVX1_1375 ( .gnd(gnd), .vdd(vdd), .A(_9831_), .Y(_10062_) );
	NAND2X1 NAND2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_9650_), .B(_9648_), .Y(_10063_) );
	OAI21X1 OAI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .B(_10035_), .C(_10063_), .Y(_10064_) );
	INVX1 INVX1_1376 ( .gnd(gnd), .vdd(vdd), .A(_10064_), .Y(_10065_) );
	NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_10062_), .B(_10065_), .Y(_10066_) );
	NAND2X1 NAND2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_10061_), .B(_10066_), .Y(_10067_) );
	INVX1 INVX1_1377 ( .gnd(gnd), .vdd(vdd), .A(_10061_), .Y(_10068_) );
	OAI21X1 OAI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_10062_), .B(_10065_), .C(_10068_), .Y(_10070_) );
	NAND3X1 NAND3X1_2149 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf1), .B(_10070_), .C(_10067_), .Y(_10071_) );
	AOI21X1 AOI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_10071_), .B(_10060_), .C(_2053_), .Y(_10072_) );
	NAND3X1 NAND3X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_10060_), .C(_10071_), .Y(_10073_) );
	NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .B(_10035_), .Y(_10074_) );
	NAND3X1 NAND3X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_9648_), .B(_9650_), .C(_10074_), .Y(_10075_) );
	NAND2X1 NAND2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_10064_), .B(_10075_), .Y(_10076_) );
	NAND2X1 NAND2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_9647_), .B(_9913__bF_buf5), .Y(_10077_) );
	OAI21X1 OAI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_9913__bF_buf4), .B(_10076_), .C(_10077_), .Y(_10078_) );
	NAND2X1 NAND2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_2042__bF_buf3), .B(_10078_), .Y(_10079_) );
	AOI21X1 AOI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_10073_), .B(_10079_), .C(_10072_), .Y(_10081_) );
	NAND3X1 NAND3X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_7453_), .B(_10032_), .C(_10043_), .Y(_10082_) );
	AOI21X1 AOI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_10043_), .B(_10032_), .C(_7453_), .Y(_10083_) );
	NAND2X1 NAND2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_10055_), .Y(_10084_) );
	OAI21X1 OAI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_10084_), .B(_10083_), .C(_10082_), .Y(_10085_) );
	AOI21X1 AOI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_10059_), .B(_10081_), .C(_10085_), .Y(_10086_) );
	OAI21X1 OAI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(divider_divuResult_2_bF_buf3), .C(_9594_), .Y(_10087_) );
	OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf0), .B(_10087_), .Y(_10088_) );
	NAND2X1 NAND2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_9591_), .B(_9598_), .Y(_10089_) );
	INVX1 INVX1_1378 ( .gnd(gnd), .vdd(vdd), .A(_9881_), .Y(_10090_) );
	OAI21X1 OAI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_9830_), .B(_10035_), .C(_9885_), .Y(_10092_) );
	AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_10092_), .B(_9840_), .Y(_10093_) );
	OAI21X1 OAI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_10090_), .B(_10093_), .C(_9843_), .Y(_10094_) );
	AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_10094_), .B(_10089_), .Y(_10095_) );
	NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_10089_), .B(_10094_), .Y(_10096_) );
	OAI21X1 OAI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_10096_), .B(_10095_), .C(divider_divuResult_1_bF_buf6), .Y(_10097_) );
	NAND3X1 NAND3X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_10088_), .C(_10097_), .Y(_10098_) );
	NAND2X1 NAND2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_10087_), .B(_9913__bF_buf3), .Y(_10099_) );
	NAND2X1 NAND2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_10089_), .B(_10094_), .Y(_10100_) );
	OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_10094_), .B(_10089_), .Y(_10101_) );
	NAND3X1 NAND3X1_2154 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf5), .B(_10100_), .C(_10101_), .Y(_10103_) );
	NAND3X1 NAND3X1_2155 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_29_), .B(_10099_), .C(_10103_), .Y(_10104_) );
	AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_10098_), .B(_10104_), .Y(_10105_) );
	OAI21X1 OAI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_9668_), .B(_10074_), .C(_9840_), .Y(_10106_) );
	NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_9881_), .B(_10106_), .Y(_10107_) );
	OAI21X1 OAI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_10090_), .B(_10093_), .C(divider_divuResult_1_bF_buf4), .Y(_10108_) );
	NAND2X1 NAND2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_9604_), .B(_9913__bF_buf2), .Y(_10109_) );
	OAI21X1 OAI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_10107_), .B(_10108_), .C(_10109_), .Y(_10110_) );
	NAND2X1 NAND2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_10110_), .Y(_10111_) );
	INVX1 INVX1_1379 ( .gnd(gnd), .vdd(vdd), .A(_10110_), .Y(_10112_) );
	NAND2X1 NAND2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_28_), .B(_10112_), .Y(_10114_) );
	AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_10114_), .B(_10111_), .Y(_10115_) );
	OAI21X1 OAI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_2240__bF_buf3), .B(_9551_), .C(divider_absoluteValue_B_flipSign_result_31_), .Y(_10116_) );
	OAI21X1 OAI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_9554_), .B(divider_divuResult_1_bF_buf3), .C(_2229__bF_buf3), .Y(_10117_) );
	INVX1 INVX1_1380 ( .gnd(gnd), .vdd(vdd), .A(_10117_), .Y(_10118_) );
	NAND2X1 NAND2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf1), .B(_10118_), .Y(_10119_) );
	NAND2X1 NAND2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_9580_), .B(_9573_), .Y(_10120_) );
	INVX1 INVX1_1381 ( .gnd(gnd), .vdd(vdd), .A(_10120_), .Y(_10121_) );
	AOI21X1 AOI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_10106_), .B(_9610_), .C(_9844_), .Y(_10122_) );
	AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_10122_), .B(_10121_), .Y(_10123_) );
	OAI21X1 OAI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_10121_), .B(_10122_), .C(divider_divuResult_1_bF_buf2), .Y(_10125_) );
	NAND3X1 NAND3X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_9570_), .B(_9572_), .C(_9913__bF_buf1), .Y(_10126_) );
	OAI21X1 OAI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_10123_), .B(_10125_), .C(_10126_), .Y(_10127_) );
	NAND2X1 NAND2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_30_), .B(_10127_), .Y(_10128_) );
	OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_10127_), .B(divider_absoluteValue_B_flipSign_result_30_), .Y(_10129_) );
	AOI22X1 AOI22X1_228 ( .gnd(gnd), .vdd(vdd), .A(_10116_), .B(_10119_), .C(_10128_), .D(_10129_), .Y(_10130_) );
	NAND3X1 NAND3X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_10115_), .B(_10105_), .C(_10130_), .Y(_10131_) );
	NAND2X1 NAND2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_10116_), .B(_10119_), .Y(_10132_) );
	NAND3X1 NAND3X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_10132_), .C(_10127_), .Y(_10133_) );
	OAI21X1 OAI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_31_), .B(_10118_), .C(_10133_), .Y(_10134_) );
	AOI21X1 AOI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_10097_), .B(_10088_), .C(_1538_), .Y(_10136_) );
	OAI21X1 OAI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10136_), .C(_10098_), .Y(_10137_) );
	AOI21X1 AOI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_10130_), .B(_10137_), .C(_10134_), .Y(_10138_) );
	OAI21X1 OAI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_10086_), .B(_10131_), .C(_10138_), .Y(_10139_) );
	NAND3X1 NAND3X1_2159 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_25_), .B(_10060_), .C(_10071_), .Y(_10140_) );
	NAND2X1 NAND2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_10060_), .B(_10071_), .Y(_10141_) );
	NAND2X1 NAND2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_2053_), .B(_10141_), .Y(_10142_) );
	INVX1 INVX1_1382 ( .gnd(gnd), .vdd(vdd), .A(_10078_), .Y(_10143_) );
	NAND2X1 NAND2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf0), .B(_10143_), .Y(_10144_) );
	NAND2X1 NAND2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_10079_), .B(_10144_), .Y(_10145_) );
	AOI21X1 AOI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_10142_), .B(_10140_), .C(_10145_), .Y(_10147_) );
	NAND2X1 NAND2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_10147_), .B(_10059_), .Y(_10148_) );
	NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .B(_10131_), .Y(_10149_) );
	AOI21X1 AOI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_10149_), .B(_10030_), .C(_10139_), .Y(_10150_) );
	NAND2X1 NAND2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_1_), .B(_1746__bF_buf5), .Y(_10151_) );
	AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .B(_10151_), .Y(_10152_) );
	NAND2X1 NAND2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_10152_), .B(divider_divuResult_1_bF_buf1), .Y(_10153_) );
	INVX1 INVX1_1383 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_1_), .Y(_10154_) );
	NAND2X1 NAND2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_10154_), .B(_9913__bF_buf0), .Y(_10155_) );
	NAND3X1 NAND3X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_1768__bF_buf3), .B(_10155_), .C(_10153_), .Y(_10156_) );
	NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_0_), .B(_1746__bF_buf4), .Y(_10158_) );
	AOI21X1 AOI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_10153_), .B(_10155_), .C(_1768__bF_buf2), .Y(_10159_) );
	OAI21X1 OAI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_10158_), .B(_10159_), .C(_10156_), .Y(_10160_) );
	XNOR2X1 XNOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_9868_), .Y(_10161_) );
	INVX1 INVX1_1384 ( .gnd(gnd), .vdd(vdd), .A(_10161_), .Y(_10162_) );
	NAND2X1 NAND2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_10162_), .B(divider_divuResult_1_bF_buf0), .Y(_10163_) );
	OAI21X1 OAI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .B(_9327_), .C(_9913__bF_buf5), .Y(_10164_) );
	NAND3X1 NAND3X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf1), .B(_10164_), .C(_10163_), .Y(_10165_) );
	NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_10161_), .B(_9913__bF_buf4), .Y(_10166_) );
	NAND2X1 NAND2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_9800_), .B(_9853_), .Y(_10167_) );
	AOI22X1 AOI22X1_229 ( .gnd(gnd), .vdd(vdd), .A(_9237_), .B(_9865_), .C(_1560__bF_buf0), .D(_10167_), .Y(_10169_) );
	OAI21X1 OAI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_10169_), .B(_10166_), .C(divider_absoluteValue_B_flipSign_result_3_bF_buf1), .Y(_10170_) );
	AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_10170_), .B(_10165_), .Y(_10171_) );
	XNOR2X1 XNOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_9864_), .B(_9334_), .Y(_10172_) );
	INVX1 INVX1_1385 ( .gnd(gnd), .vdd(vdd), .A(_10172_), .Y(_10173_) );
	NAND3X1 NAND3X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf3), .B(_10173_), .C(_10167_), .Y(_10174_) );
	OAI21X1 OAI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_9030_), .B(_9325__bF_buf3), .C(_9330_), .Y(_10175_) );
	INVX1 INVX1_1386 ( .gnd(gnd), .vdd(vdd), .A(_10175_), .Y(_10176_) );
	NAND2X1 NAND2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_9913__bF_buf3), .Y(_10177_) );
	NAND3X1 NAND3X1_2163 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_2_bF_buf1), .B(_10174_), .C(_10177_), .Y(_10178_) );
	NAND2X1 NAND2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_10175_), .B(_9913__bF_buf2), .Y(_10180_) );
	NAND3X1 NAND3X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf2), .B(_10172_), .C(_10167_), .Y(_10181_) );
	NAND3X1 NAND3X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_2547__bF_buf3), .B(_10181_), .C(_10180_), .Y(_10182_) );
	NAND2X1 NAND2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_10178_), .B(_10182_), .Y(_10183_) );
	NAND3X1 NAND3X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_10183_), .B(_10160_), .C(_10171_), .Y(_10184_) );
	INVX1 INVX1_1387 ( .gnd(gnd), .vdd(vdd), .A(_10165_), .Y(_10185_) );
	AOI21X1 AOI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_10180_), .B(_10181_), .C(divider_absoluteValue_B_flipSign_result_2_bF_buf0), .Y(_10186_) );
	AOI21X1 AOI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_10170_), .B(_10186_), .C(_10185_), .Y(_10187_) );
	NAND2X1 NAND2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_9913__bF_buf1), .Y(_10188_) );
	NAND2X1 NAND2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_9353_), .Y(_10189_) );
	NAND2X1 NAND2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_9393_), .B(_9338_), .Y(_10191_) );
	AOI22X1 AOI22X1_230 ( .gnd(gnd), .vdd(vdd), .A(_9359_), .B(_9362_), .C(_9404_), .D(_10191_), .Y(_10192_) );
	OAI21X1 OAI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_9408_), .B(_10192_), .C(_10189_), .Y(_10193_) );
	INVX1 INVX1_1388 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .Y(_10194_) );
	INVX1 INVX1_1389 ( .gnd(gnd), .vdd(vdd), .A(_9408_), .Y(_10195_) );
	NAND2X1 NAND2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_9359_), .B(_9362_), .Y(_10196_) );
	NAND2X1 NAND2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_10191_), .Y(_10197_) );
	NAND2X1 NAND2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_10196_), .B(_10197_), .Y(_10198_) );
	NAND3X1 NAND3X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_10194_), .B(_10195_), .C(_10198_), .Y(_10199_) );
	NAND2X1 NAND2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_10193_), .B(_10199_), .Y(_10200_) );
	NAND3X1 NAND3X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf1), .B(_10200_), .C(_10167_), .Y(_10202_) );
	NAND3X1 NAND3X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_4714__bF_buf0), .B(_10202_), .C(_10188_), .Y(_10203_) );
	INVX1 INVX1_1390 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .Y(_10204_) );
	NAND2X1 NAND2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_10204_), .B(_9913__bF_buf0), .Y(_10205_) );
	NAND3X1 NAND3X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .B(_10195_), .C(_10198_), .Y(_10206_) );
	OAI21X1 OAI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_9408_), .B(_10192_), .C(_10194_), .Y(_10207_) );
	NAND2X1 NAND2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_10207_), .B(_10206_), .Y(_10208_) );
	NAND3X1 NAND3X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf0), .B(_10208_), .C(_10167_), .Y(_10209_) );
	NAND3X1 NAND3X1_2172 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_7_bF_buf0), .B(_10209_), .C(_10205_), .Y(_10210_) );
	NAND2X1 NAND2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_10203_), .B(_10210_), .Y(_10211_) );
	NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_10196_), .B(_10197_), .Y(_10213_) );
	NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_10192_), .B(_10213_), .Y(_10214_) );
	INVX1 INVX1_1391 ( .gnd(gnd), .vdd(vdd), .A(_10214_), .Y(_10215_) );
	NAND3X1 NAND3X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf3), .B(_10215_), .C(_10167_), .Y(_10216_) );
	OAI21X1 OAI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf2), .B(_9354_), .C(_9358_), .Y(_10217_) );
	NAND2X1 NAND2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_10217_), .B(_9913__bF_buf5), .Y(_10218_) );
	NAND3X1 NAND3X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_4999__bF_buf1), .B(_10216_), .C(_10218_), .Y(_10219_) );
	NAND3X1 NAND3X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf2), .B(_10214_), .C(_10167_), .Y(_10220_) );
	INVX1 INVX1_1392 ( .gnd(gnd), .vdd(vdd), .A(_10217_), .Y(_10221_) );
	NAND2X1 NAND2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_10221_), .B(_9913__bF_buf4), .Y(_10222_) );
	NAND3X1 NAND3X1_2176 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf2), .B(_10220_), .C(_10222_), .Y(_10224_) );
	NAND2X1 NAND2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_10224_), .B(_10219_), .Y(_10225_) );
	NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_10211_), .B(_10225_), .Y(_10226_) );
	NAND2X1 NAND2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_9391_), .B(_9913__bF_buf3), .Y(_10227_) );
	NAND2X1 NAND2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_9392_), .Y(_10228_) );
	INVX1 INVX1_1393 ( .gnd(gnd), .vdd(vdd), .A(_9338_), .Y(_10229_) );
	INVX1 INVX1_1394 ( .gnd(gnd), .vdd(vdd), .A(_9402_), .Y(_10230_) );
	NAND2X1 NAND2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_2470__bF_buf0), .B(_10230_), .Y(_10231_) );
	AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_9381_), .B(_9378_), .Y(_10232_) );
	OAI21X1 OAI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_10232_), .B(_10229_), .C(_10231_), .Y(_10233_) );
	XNOR2X1 XNOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_10233_), .B(_10228_), .Y(_10235_) );
	NAND3X1 NAND3X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf1), .B(_10235_), .C(_10167_), .Y(_10236_) );
	NAND3X1 NAND3X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_4100__bF_buf0), .B(_10236_), .C(_10227_), .Y(_10237_) );
	NAND2X1 NAND2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_9913__bF_buf2), .Y(_10238_) );
	XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_10233_), .B(_10228_), .Y(_10239_) );
	NAND3X1 NAND3X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf0), .B(_10239_), .C(_10167_), .Y(_10240_) );
	NAND3X1 NAND3X1_2180 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_5_bF_buf0), .B(_10240_), .C(_10238_), .Y(_10241_) );
	NAND2X1 NAND2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_10237_), .B(_10241_), .Y(_10242_) );
	XNOR2X1 XNOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_9338_), .B(_10232_), .Y(_10243_) );
	INVX1 INVX1_1395 ( .gnd(gnd), .vdd(vdd), .A(_10243_), .Y(_10244_) );
	NAND3X1 NAND3X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf3), .B(_10244_), .C(_10167_), .Y(_10246_) );
	NAND2X1 NAND2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_9402_), .B(_9913__bF_buf1), .Y(_10247_) );
	NAND3X1 NAND3X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_10246_), .C(_10247_), .Y(_10248_) );
	NAND2X1 NAND2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_10230_), .B(_9913__bF_buf0), .Y(_10249_) );
	NAND3X1 NAND3X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf2), .B(_10243_), .C(_10167_), .Y(_10250_) );
	NAND3X1 NAND3X1_2184 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_4_bF_buf6), .B(_10250_), .C(_10249_), .Y(_10251_) );
	NAND2X1 NAND2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_10248_), .B(_10251_), .Y(_10252_) );
	NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_10242_), .B(_10252_), .Y(_10253_) );
	NAND2X1 NAND2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_10226_), .B(_10253_), .Y(_10254_) );
	AOI21X1 AOI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_10184_), .B(_10187_), .C(_10254_), .Y(_10255_) );
	OAI21X1 OAI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_10221_), .B(divider_divuResult_1_bF_buf6), .C(_10216_), .Y(_10257_) );
	OAI21X1 OAI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf1), .B(_10257_), .C(_10203_), .Y(_10258_) );
	OAI21X1 OAI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_10248_), .B(_10242_), .C(_10237_), .Y(_10259_) );
	AOI22X1 AOI22X1_231 ( .gnd(gnd), .vdd(vdd), .A(_10210_), .B(_10258_), .C(_10226_), .D(_10259_), .Y(_10260_) );
	INVX1 INVX1_1396 ( .gnd(gnd), .vdd(vdd), .A(_10260_), .Y(_10261_) );
	NAND2X1 NAND2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_9544_), .B(_9913__bF_buf5), .Y(_10262_) );
	INVX1 INVX1_1397 ( .gnd(gnd), .vdd(vdd), .A(_9546_), .Y(_10263_) );
	NAND2X1 NAND2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_9441_), .Y(_10264_) );
	INVX1 INVX1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9543_), .Y(_10265_) );
	INVX1 INVX1_1399 ( .gnd(gnd), .vdd(vdd), .A(_9467_), .Y(_10266_) );
	INVX1 INVX1_1400 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .Y(_10268_) );
	OAI21X1 OAI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9872_), .C(_9516_), .Y(_10269_) );
	AOI21X1 AOI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_10269_), .B(_10268_), .C(_10266_), .Y(_10270_) );
	OAI21X1 OAI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_10265_), .B(_10270_), .C(_10264_), .Y(_10271_) );
	NAND3X1 NAND3X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_9534_), .B(_10263_), .C(_10271_), .Y(_10272_) );
	INVX1 INVX1_1401 ( .gnd(gnd), .vdd(vdd), .A(_9534_), .Y(_10273_) );
	INVX1 INVX1_1402 ( .gnd(gnd), .vdd(vdd), .A(_10264_), .Y(_10274_) );
	INVX1 INVX1_1403 ( .gnd(gnd), .vdd(vdd), .A(_9541_), .Y(_10275_) );
	OAI21X1 OAI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf0), .B(_9538_), .C(_10275_), .Y(_10276_) );
	OAI21X1 OAI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_9874_), .B(_9412_), .C(_10268_), .Y(_10277_) );
	AOI22X1 AOI22X1_232 ( .gnd(gnd), .vdd(vdd), .A(_9540_), .B(_10276_), .C(_9467_), .D(_10277_), .Y(_10279_) );
	OAI21X1 OAI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_10274_), .B(_10279_), .C(_10263_), .Y(_10280_) );
	NAND2X1 NAND2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_10273_), .B(_10280_), .Y(_10281_) );
	NAND3X1 NAND3X1_2186 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf5), .B(_10272_), .C(_10281_), .Y(_10282_) );
	NAND3X1 NAND3X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_1944__bF_buf1), .B(_10262_), .C(_10282_), .Y(_10283_) );
	INVX1 INVX1_1404 ( .gnd(gnd), .vdd(vdd), .A(_9544_), .Y(_10284_) );
	NAND2X1 NAND2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_10284_), .B(_9913__bF_buf4), .Y(_10285_) );
	NAND2X1 NAND2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_9534_), .B(_10280_), .Y(_10286_) );
	NAND3X1 NAND3X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_10273_), .B(_10263_), .C(_10271_), .Y(_10287_) );
	NAND3X1 NAND3X1_2189 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf4), .B(_10287_), .C(_10286_), .Y(_10288_) );
	NAND3X1 NAND3X1_2190 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_15_bF_buf1), .B(_10285_), .C(_10288_), .Y(_10290_) );
	AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_10283_), .B(_10290_), .Y(_10291_) );
	NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_10274_), .B(_10279_), .Y(_10292_) );
	AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_10279_), .B(_10274_), .Y(_10293_) );
	OAI21X1 OAI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10293_), .C(divider_divuResult_1_bF_buf3), .Y(_10294_) );
	NAND2X1 NAND2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_9440_), .B(_9913__bF_buf3), .Y(_10295_) );
	NAND3X1 NAND3X1_2191 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf4), .B(_10295_), .C(_10294_), .Y(_10296_) );
	NAND2X1 NAND2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_10274_), .B(_10279_), .Y(_10297_) );
	NAND3X1 NAND3X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_10271_), .B(_10297_), .C(divider_divuResult_1_bF_buf2), .Y(_10298_) );
	INVX1 INVX1_1405 ( .gnd(gnd), .vdd(vdd), .A(_9440_), .Y(_10299_) );
	NAND2X1 NAND2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_10299_), .B(_9913__bF_buf2), .Y(_10301_) );
	NAND3X1 NAND3X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf4), .B(_10301_), .C(_10298_), .Y(_10302_) );
	NAND2X1 NAND2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_10302_), .B(_10296_), .Y(_10303_) );
	OAI21X1 OAI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_9455_), .B(_9456_), .C(_9913__bF_buf1), .Y(_10304_) );
	NAND2X1 NAND2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_9452_), .B(_9457_), .Y(_10305_) );
	INVX1 INVX1_1406 ( .gnd(gnd), .vdd(vdd), .A(_10305_), .Y(_10306_) );
	NAND2X1 NAND2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_9462_), .B(_9466_), .Y(_10307_) );
	NAND2X1 NAND2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_10307_), .B(_10277_), .Y(_10308_) );
	AOI21X1 AOI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_10308_), .B(_10275_), .C(_10306_), .Y(_10309_) );
	AOI22X1 AOI22X1_233 ( .gnd(gnd), .vdd(vdd), .A(_9462_), .B(_9466_), .C(_10268_), .D(_10269_), .Y(_10310_) );
	NOR3X1 NOR3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_10305_), .B(_9541_), .C(_10310_), .Y(_10312_) );
	OAI21X1 OAI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_10309_), .B(_10312_), .C(divider_divuResult_1_bF_buf1), .Y(_10313_) );
	NAND3X1 NAND3X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_1494__bF_buf0), .B(_10304_), .C(_10313_), .Y(_10314_) );
	INVX1 INVX1_1407 ( .gnd(gnd), .vdd(vdd), .A(_9538_), .Y(_10315_) );
	NAND2X1 NAND2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_10315_), .B(_9913__bF_buf0), .Y(_10316_) );
	NOR3X1 NOR3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_10306_), .B(_9541_), .C(_10310_), .Y(_10317_) );
	AOI21X1 AOI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_10308_), .B(_10275_), .C(_10305_), .Y(_10318_) );
	OAI21X1 OAI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_10317_), .B(_10318_), .C(divider_divuResult_1_bF_buf0), .Y(_10319_) );
	NAND3X1 NAND3X1_2195 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf5), .B(_10316_), .C(_10319_), .Y(_10320_) );
	NAND2X1 NAND2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_10314_), .B(_10320_), .Y(_10321_) );
	XNOR2X1 XNOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_10277_), .B(_10307_), .Y(_10323_) );
	NAND3X1 NAND3X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf1), .B(_10323_), .C(_10167_), .Y(_10324_) );
	NAND2X1 NAND2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_9461_), .Y(_10325_) );
	NAND2X1 NAND2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_10325_), .B(_9913__bF_buf5), .Y(_10326_) );
	NAND3X1 NAND3X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_1484__bF_buf4), .B(_10324_), .C(_10326_), .Y(_10327_) );
	NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_10307_), .B(_10277_), .Y(_10328_) );
	NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_10310_), .B(_10328_), .Y(_10329_) );
	NAND3X1 NAND3X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf0), .B(_10167_), .C(_10329_), .Y(_10330_) );
	INVX1 INVX1_1408 ( .gnd(gnd), .vdd(vdd), .A(_10325_), .Y(_10331_) );
	NAND2X1 NAND2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_10331_), .B(_9913__bF_buf4), .Y(_10332_) );
	NAND3X1 NAND3X1_2199 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_12_bF_buf5), .B(_10330_), .C(_10332_), .Y(_10334_) );
	NAND2X1 NAND2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_10327_), .B(_10334_), .Y(_10335_) );
	NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_10335_), .B(_10321_), .Y(_10336_) );
	NAND3X1 NAND3X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_10303_), .B(_10336_), .C(_10291_), .Y(_10337_) );
	OAI21X1 OAI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_9483_), .C(_9913__bF_buf3), .Y(_10338_) );
	NAND2X1 NAND2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_9481_), .B(_9484_), .Y(_10339_) );
	INVX1 INVX1_1409 ( .gnd(gnd), .vdd(vdd), .A(_10339_), .Y(_10340_) );
	INVX1 INVX1_1410 ( .gnd(gnd), .vdd(vdd), .A(_9526_), .Y(_10341_) );
	INVX1 INVX1_1411 ( .gnd(gnd), .vdd(vdd), .A(_9515_), .Y(_10342_) );
	OAI21X1 OAI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_10342_), .B(_9412_), .C(_9532_), .Y(_10343_) );
	NAND2X1 NAND2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_9521_), .B(_10343_), .Y(_10345_) );
	AOI21X1 AOI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_10345_), .B(_10341_), .C(_10340_), .Y(_10346_) );
	NAND3X1 NAND3X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_10340_), .B(_10341_), .C(_10345_), .Y(_10347_) );
	INVX1 INVX1_1412 ( .gnd(gnd), .vdd(vdd), .A(_10347_), .Y(_10348_) );
	OAI21X1 OAI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_10346_), .B(_10348_), .C(divider_divuResult_1_bF_buf6), .Y(_10349_) );
	NAND3X1 NAND3X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_1265__bF_buf2), .B(_10338_), .C(_10349_), .Y(_10350_) );
	AOI21X1 AOI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_9469_), .B(_9480_), .C(divider_divuResult_1_bF_buf5), .Y(_10351_) );
	AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_10343_), .B(_9521_), .Y(_10352_) );
	OAI21X1 OAI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_9526_), .B(_10352_), .C(_10339_), .Y(_10353_) );
	AOI21X1 AOI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_10353_), .B(_10347_), .C(_9913__bF_buf2), .Y(_10354_) );
	OAI21X1 OAI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_10351_), .B(_10354_), .C(divider_absoluteValue_B_flipSign_result_11_bF_buf3), .Y(_10356_) );
	AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_10356_), .B(_10350_), .Y(_10357_) );
	NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_9521_), .B(_10343_), .Y(_10358_) );
	OAI21X1 OAI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_10352_), .B(_10358_), .C(divider_divuResult_1_bF_buf4), .Y(_10359_) );
	NAND2X1 NAND2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_9525_), .B(_9913__bF_buf1), .Y(_10360_) );
	NAND3X1 NAND3X1_2203 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_10_bF_buf1), .B(_10360_), .C(_10359_), .Y(_10361_) );
	NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_10358_), .B(_10352_), .Y(_10362_) );
	NAND2X1 NAND2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_10362_), .B(divider_divuResult_1_bF_buf3), .Y(_10363_) );
	NAND3X1 NAND3X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_9488_), .B(_9489_), .C(_9913__bF_buf0), .Y(_10364_) );
	NAND3X1 NAND3X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_10678__bF_buf5), .B(_10363_), .C(_10364_), .Y(_10365_) );
	NAND2X1 NAND2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_10361_), .B(_10365_), .Y(_10367_) );
	NAND3X1 NAND3X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_9506_), .B(_9511_), .C(_9913__bF_buf5), .Y(_10368_) );
	INVX1 INVX1_1413 ( .gnd(gnd), .vdd(vdd), .A(_9529_), .Y(_10369_) );
	INVX1 INVX1_1414 ( .gnd(gnd), .vdd(vdd), .A(_9528_), .Y(_10370_) );
	NAND2X1 NAND2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_9504_), .B(_9501_), .Y(_10371_) );
	INVX1 INVX1_1415 ( .gnd(gnd), .vdd(vdd), .A(_10371_), .Y(_10372_) );
	OAI21X1 OAI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_10372_), .B(_9412_), .C(_10370_), .Y(_10373_) );
	NAND3X1 NAND3X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_10369_), .B(_9530_), .C(_10373_), .Y(_10374_) );
	NAND2X1 NAND2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_9530_), .B(_10369_), .Y(_10375_) );
	OAI21X1 OAI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_9872_), .C(_10371_), .Y(_10376_) );
	NAND3X1 NAND3X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_10370_), .B(_10375_), .C(_10376_), .Y(_10378_) );
	NAND2X1 NAND2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_10378_), .B(_10374_), .Y(_10379_) );
	NAND3X1 NAND3X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_1560__bF_buf3), .B(_10379_), .C(_10167_), .Y(_10380_) );
	NAND3X1 NAND3X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_8971__bF_buf0), .B(_10380_), .C(_10368_), .Y(_10381_) );
	NAND2X1 NAND2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_9512_), .B(_9913__bF_buf4), .Y(_10382_) );
	INVX1 INVX1_1416 ( .gnd(gnd), .vdd(vdd), .A(_10379_), .Y(_10383_) );
	NAND2X1 NAND2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf2), .B(_10383_), .Y(_10384_) );
	NAND3X1 NAND3X1_2211 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_9_bF_buf2), .B(_10382_), .C(_10384_), .Y(_10385_) );
	NAND2X1 NAND2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_10385_), .Y(_10386_) );
	NAND2X1 NAND2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_10372_), .B(_9412_), .Y(_10387_) );
	NAND2X1 NAND2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_10376_), .B(_10387_), .Y(_10389_) );
	NAND2X1 NAND2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_10389_), .B(divider_divuResult_1_bF_buf1), .Y(_10390_) );
	OAI21X1 OAI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_9325__bF_buf1), .B(_9497_), .C(_9500_), .Y(_10391_) );
	NAND2X1 NAND2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_10391_), .B(_9913__bF_buf3), .Y(_10392_) );
	NAND3X1 NAND3X1_2212 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf3), .B(_10392_), .C(_10390_), .Y(_10393_) );
	NAND3X1 NAND3X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_9499_), .B(_9500_), .C(_9913__bF_buf2), .Y(_10394_) );
	INVX1 INVX1_1417 ( .gnd(gnd), .vdd(vdd), .A(_10389_), .Y(_10395_) );
	NAND2X1 NAND2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_10395_), .B(divider_divuResult_1_bF_buf0), .Y(_10396_) );
	NAND3X1 NAND3X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_7204__bF_buf0), .B(_10396_), .C(_10394_), .Y(_10397_) );
	AOI21X1 AOI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_10393_), .B(_10397_), .C(_10386_), .Y(_10398_) );
	NAND3X1 NAND3X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_10357_), .B(_10367_), .C(_10398_), .Y(_10400_) );
	NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_10400_), .B(_10337_), .Y(_10401_) );
	OAI21X1 OAI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(_10261_), .C(_10401_), .Y(_10402_) );
	NAND3X1 NAND3X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_10283_), .B(_10290_), .C(_10303_), .Y(_10403_) );
	INVX1 INVX1_1418 ( .gnd(gnd), .vdd(vdd), .A(_10336_), .Y(_10404_) );
	NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_10403_), .B(_10404_), .Y(_10405_) );
	NAND3X1 NAND3X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_10350_), .B(_10356_), .C(_10367_), .Y(_10406_) );
	OAI21X1 OAI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_9913__bF_buf1), .B(_10395_), .C(_10392_), .Y(_10407_) );
	OAI21X1 OAI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf2), .B(_10407_), .C(_10381_), .Y(_10408_) );
	NAND2X1 NAND2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_10385_), .B(_10408_), .Y(_10409_) );
	INVX1 INVX1_1419 ( .gnd(gnd), .vdd(vdd), .A(_10350_), .Y(_10411_) );
	AOI21X1 AOI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_10364_), .B(_10363_), .C(divider_absoluteValue_B_flipSign_result_10_bF_buf0), .Y(_10412_) );
	AOI21X1 AOI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_10412_), .B(_10356_), .C(_10411_), .Y(_10413_) );
	OAI21X1 OAI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_10409_), .B(_10406_), .C(_10413_), .Y(_10414_) );
	OAI21X1 OAI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_10315_), .B(divider_divuResult_1_bF_buf6), .C(_10313_), .Y(_10415_) );
	OAI21X1 OAI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_13_bF_buf4), .B(_10415_), .C(_10327_), .Y(_10416_) );
	NAND2X1 NAND2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_10320_), .B(_10416_), .Y(_10417_) );
	AOI21X1 AOI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_10288_), .B(_10285_), .C(divider_absoluteValue_B_flipSign_result_15_bF_buf0), .Y(_10418_) );
	NAND3X1 NAND3X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_1505__bF_buf3), .B(_10295_), .C(_10294_), .Y(_10419_) );
	INVX1 INVX1_1420 ( .gnd(gnd), .vdd(vdd), .A(_10419_), .Y(_10420_) );
	AOI21X1 AOI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .B(_10290_), .C(_10418_), .Y(_10422_) );
	OAI21X1 OAI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_10417_), .B(_10403_), .C(_10422_), .Y(_10423_) );
	AOI21X1 AOI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_10405_), .B(_10414_), .C(_10423_), .Y(_10424_) );
	NAND2X1 NAND2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_10424_), .B(_10402_), .Y(_10425_) );
	NAND2X1 NAND2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_9939_), .B(_9942_), .Y(_10426_) );
	NAND3X1 NAND3X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_10022_), .B(_10023_), .C(_10426_), .Y(_10427_) );
	INVX1 INVX1_1421 ( .gnd(gnd), .vdd(vdd), .A(_10005_), .Y(_10428_) );
	INVX1 INVX1_1422 ( .gnd(gnd), .vdd(vdd), .A(_10007_), .Y(_10429_) );
	NAND3X1 NAND3X1_2220 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf0), .B(_10429_), .C(_10428_), .Y(_10430_) );
	NAND2X1 NAND2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_10008_), .B(_10430_), .Y(_10431_) );
	NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_10431_), .B(_10011_), .Y(_10433_) );
	NAND2X1 NAND2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_9993_), .B(_10433_), .Y(_10434_) );
	NOR3X1 NOR3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_9962_), .B(_10427_), .C(_10434_), .Y(_10435_) );
	NAND3X1 NAND3X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_10425_), .B(_10435_), .C(_10149_), .Y(_10436_) );
	NAND2X1 NAND2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_10436_), .B(_10150_), .Y(divider_divuResult_0_) );
	INVX1 INVX1_1423 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_0_), .Y(_10437_) );
	NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf2), .B(_10437_), .Y(_10438_) );
	OAI21X1 OAI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_10158_), .B(_10438_), .C(divider_divuResult_0_bF_buf6), .Y(_10439_) );
	OAI21X1 OAI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_10437_), .B(divider_divuResult_0_bF_buf5), .C(_10439_), .Y(divider_flipSign_rem_operand_0_) );
	INVX1 INVX1_1424 ( .gnd(gnd), .vdd(vdd), .A(_10152_), .Y(_10440_) );
	NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_10440_), .B(_9913__bF_buf0), .Y(_10442_) );
	NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(divider_aOp_abs_1_), .B(divider_divuResult_1_bF_buf5), .Y(_10443_) );
	OAI21X1 OAI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_10442_), .B(_10443_), .C(divider_absoluteValue_B_flipSign_result_1_bF_buf7), .Y(_10444_) );
	NAND2X1 NAND2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_10156_), .B(_10444_), .Y(_10445_) );
	XNOR2X1 XNOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_10445_), .B(_10158_), .Y(_10446_) );
	AOI21X1 AOI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_10153_), .B(_10155_), .C(divider_divuResult_0_bF_buf4), .Y(_10447_) );
	AOI21X1 AOI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf3), .B(_10446_), .C(_10447_), .Y(divider_flipSign_rem_operand_1_) );
	XNOR2X1 XNOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_10160_), .B(_10183_), .Y(_10448_) );
	AOI21X1 AOI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_10174_), .B(_10177_), .C(divider_divuResult_0_bF_buf2), .Y(_10449_) );
	AOI21X1 AOI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf1), .B(_10448_), .C(_10449_), .Y(divider_flipSign_rem_operand_2_) );
	AOI21X1 AOI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_10160_), .B(_10183_), .C(_10186_), .Y(_10451_) );
	XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_10451_), .B(_10171_), .Y(_10452_) );
	AOI21X1 AOI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_10163_), .B(_10164_), .C(divider_divuResult_0_bF_buf0), .Y(_10453_) );
	AOI21X1 AOI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf6), .B(_10452_), .C(_10453_), .Y(divider_flipSign_rem_operand_3_) );
	NOR3X1 NOR3X1_102 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_1_bF_buf6), .B(_10442_), .C(_10443_), .Y(_10454_) );
	INVX1 INVX1_1425 ( .gnd(gnd), .vdd(vdd), .A(_10158_), .Y(_10455_) );
	AOI21X1 AOI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_10455_), .B(_10444_), .C(_10454_), .Y(_10456_) );
	NAND3X1 NAND3X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_10165_), .B(_10170_), .C(_10183_), .Y(_10457_) );
	OAI21X1 OAI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_10456_), .B(_10457_), .C(_10187_), .Y(_10458_) );
	XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_10458_), .B(_10252_), .Y(_10459_) );
	AOI21X1 AOI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_10246_), .B(_10247_), .C(divider_divuResult_0_bF_buf5), .Y(_10461_) );
	AOI21X1 AOI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf4), .B(_10459_), .C(_10461_), .Y(divider_flipSign_rem_operand_4_) );
	INVX1 INVX1_1426 ( .gnd(gnd), .vdd(vdd), .A(_10458_), .Y(_10462_) );
	OAI21X1 OAI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_10252_), .B(_10462_), .C(_10248_), .Y(_10463_) );
	XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_10463_), .B(_10242_), .Y(_10464_) );
	AOI21X1 AOI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_10227_), .B(_10236_), .C(divider_divuResult_0_bF_buf3), .Y(_10465_) );
	AOI21X1 AOI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf2), .B(_10464_), .C(_10465_), .Y(divider_flipSign_rem_operand_5_) );
	INVX1 INVX1_1427 ( .gnd(gnd), .vdd(vdd), .A(_10225_), .Y(_10466_) );
	INVX1 INVX1_1428 ( .gnd(gnd), .vdd(vdd), .A(_10253_), .Y(_10467_) );
	INVX1 INVX1_1429 ( .gnd(gnd), .vdd(vdd), .A(_10259_), .Y(_10468_) );
	OAI21X1 OAI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_10467_), .B(_10462_), .C(_10468_), .Y(_10470_) );
	XNOR2X1 XNOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_10470_), .B(_10466_), .Y(_10471_) );
	MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_10471_), .B(_10257_), .S(divider_divuResult_0_bF_buf1), .Y(divider_flipSign_rem_operand_6_) );
	OAI21X1 OAI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(divider_divuResult_1_bF_buf4), .C(_10209_), .Y(_10472_) );
	INVX1 INVX1_1430 ( .gnd(gnd), .vdd(vdd), .A(_10472_), .Y(_10473_) );
	NAND2X1 NAND2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_10466_), .B(_10470_), .Y(_10474_) );
	OAI21X1 OAI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_6_bF_buf0), .B(_10257_), .C(_10474_), .Y(_10475_) );
	AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_10475_), .B(_10211_), .Y(_10476_) );
	NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_10211_), .B(_10475_), .Y(_10477_) );
	OAI21X1 OAI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_10476_), .B(_10477_), .C(divider_divuResult_0_bF_buf0), .Y(_10478_) );
	OAI21X1 OAI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_10473_), .B(divider_divuResult_0_bF_buf6), .C(_10478_), .Y(divider_flipSign_rem_operand_7_) );
	NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_10261_), .B(_10255_), .Y(_10480_) );
	NAND2X1 NAND2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_10393_), .B(_10397_), .Y(_10481_) );
	XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_10480_), .B(_10481_), .Y(_10482_) );
	MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_10482_), .B(_10407_), .S(divider_divuResult_0_bF_buf5), .Y(divider_flipSign_rem_operand_8_) );
	OAI21X1 OAI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_10261_), .B(_10255_), .C(_10481_), .Y(_10483_) );
	OAI21X1 OAI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_8_bF_buf1), .B(_10407_), .C(_10483_), .Y(_10484_) );
	XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_10484_), .B(_10386_), .Y(_10485_) );
	AOI21X1 AOI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_10368_), .B(_10380_), .C(divider_divuResult_0_bF_buf4), .Y(_10486_) );
	AOI21X1 AOI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf3), .B(_10485_), .C(_10486_), .Y(divider_flipSign_rem_operand_9_) );
	NAND3X1 NAND3X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_10381_), .B(_10385_), .C(_10481_), .Y(_10488_) );
	OAI21X1 OAI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_10488_), .B(_10480_), .C(_10409_), .Y(_10489_) );
	XNOR2X1 XNOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_10489_), .B(_10367_), .Y(_10490_) );
	AOI21X1 AOI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_10359_), .B(_10360_), .C(divider_divuResult_0_bF_buf2), .Y(_10491_) );
	AOI21X1 AOI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf1), .B(_10490_), .C(_10491_), .Y(divider_flipSign_rem_operand_10_) );
	NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_10351_), .B(_10354_), .Y(_10492_) );
	INVX1 INVX1_1431 ( .gnd(gnd), .vdd(vdd), .A(_10492_), .Y(_10493_) );
	INVX1 INVX1_1432 ( .gnd(gnd), .vdd(vdd), .A(_10412_), .Y(_10494_) );
	NAND2X1 NAND2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_10367_), .B(_10489_), .Y(_10495_) );
	NAND2X1 NAND2X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_10494_), .B(_10495_), .Y(_10496_) );
	NAND2X1 NAND2X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_10357_), .B(_10496_), .Y(_10498_) );
	OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_10496_), .B(_10357_), .Y(_10499_) );
	NAND3X1 NAND3X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_10498_), .B(_10499_), .C(divider_divuResult_0_bF_buf0), .Y(_10500_) );
	OAI21X1 OAI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_10493_), .B(divider_divuResult_0_bF_buf6), .C(_10500_), .Y(divider_flipSign_rem_operand_11_) );
	INVX1 INVX1_1433 ( .gnd(gnd), .vdd(vdd), .A(_10335_), .Y(_10501_) );
	INVX1 INVX1_1434 ( .gnd(gnd), .vdd(vdd), .A(_10414_), .Y(_10502_) );
	OAI21X1 OAI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_10400_), .B(_10480_), .C(_10502_), .Y(_10503_) );
	XNOR2X1 XNOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_10503_), .B(_10501_), .Y(_10504_) );
	AOI21X1 AOI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_10324_), .B(_10326_), .C(divider_divuResult_0_bF_buf5), .Y(_10505_) );
	AOI21X1 AOI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf4), .B(_10504_), .C(_10505_), .Y(divider_flipSign_rem_operand_12_) );
	NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_10400_), .B(_10480_), .Y(_10507_) );
	OAI21X1 OAI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_10414_), .B(_10507_), .C(_10501_), .Y(_10508_) );
	NAND2X1 NAND2X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_10327_), .B(_10508_), .Y(_10509_) );
	AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_10509_), .B(_10321_), .Y(_10510_) );
	NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_10321_), .B(_10509_), .Y(_10511_) );
	OAI21X1 OAI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_10511_), .B(_10510_), .C(divider_divuResult_0_bF_buf3), .Y(_10512_) );
	OAI21X1 OAI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_10415_), .B(divider_divuResult_0_bF_buf2), .C(_10512_), .Y(divider_flipSign_rem_operand_13_) );
	OAI21X1 OAI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_10299_), .B(divider_divuResult_1_bF_buf3), .C(_10294_), .Y(_10513_) );
	INVX1 INVX1_1435 ( .gnd(gnd), .vdd(vdd), .A(_10417_), .Y(_10514_) );
	AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_10503_), .B(_10336_), .Y(_10515_) );
	OAI21X1 OAI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_10514_), .B(_10515_), .C(_10303_), .Y(_10517_) );
	NAND3X1 NAND3X1_2225 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_14_bF_buf3), .B(_10301_), .C(_10298_), .Y(_10518_) );
	NAND2X1 NAND2X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_10518_), .B(_10419_), .Y(_10519_) );
	OAI21X1 OAI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_10414_), .B(_10507_), .C(_10336_), .Y(_10520_) );
	NAND3X1 NAND3X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .B(_10417_), .C(_10520_), .Y(_10521_) );
	NAND3X1 NAND3X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_10517_), .B(_10521_), .C(divider_divuResult_0_bF_buf1), .Y(_10522_) );
	OAI21X1 OAI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_10513_), .B(divider_divuResult_0_bF_buf0), .C(_10522_), .Y(divider_flipSign_rem_operand_14_) );
	OAI21X1 OAI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_10284_), .B(divider_divuResult_1_bF_buf2), .C(_10282_), .Y(_10523_) );
	INVX1 INVX1_1436 ( .gnd(gnd), .vdd(vdd), .A(_10291_), .Y(_10524_) );
	NAND3X1 NAND3X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_10524_), .B(_10419_), .C(_10517_), .Y(_10525_) );
	AOI21X1 AOI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_10520_), .B(_10417_), .C(_10519_), .Y(_10527_) );
	OAI21X1 OAI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_10420_), .B(_10527_), .C(_10291_), .Y(_10528_) );
	NAND3X1 NAND3X1_2229 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf6), .B(_10525_), .C(_10528_), .Y(_10529_) );
	OAI21X1 OAI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_10523_), .B(divider_divuResult_0_bF_buf5), .C(_10529_), .Y(divider_flipSign_rem_operand_15_) );
	OAI21X1 OAI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_10004_), .B(divider_divuResult_1_bF_buf1), .C(_10429_), .Y(_10530_) );
	INVX1 INVX1_1437 ( .gnd(gnd), .vdd(vdd), .A(_10530_), .Y(_10531_) );
	NAND3X1 NAND3X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_10008_), .B(_10430_), .C(_10425_), .Y(_10532_) );
	NAND3X1 NAND3X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_10424_), .B(_10431_), .C(_10402_), .Y(_10533_) );
	NAND3X1 NAND3X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_10532_), .B(_10533_), .C(divider_divuResult_0_bF_buf4), .Y(_10534_) );
	OAI21X1 OAI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_10531_), .B(divider_divuResult_0_bF_buf3), .C(_10534_), .Y(divider_flipSign_rem_operand_16_) );
	INVX1 INVX1_1438 ( .gnd(gnd), .vdd(vdd), .A(_10001_), .Y(_10536_) );
	OAI21X1 OAI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_16_bF_buf5), .B(_10531_), .C(_10532_), .Y(_10537_) );
	XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_10537_), .B(_10011_), .Y(_10538_) );
	MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_10538_), .B(_10536_), .S(divider_divuResult_0_bF_buf2), .Y(divider_flipSign_rem_operand_17_) );
	AOI21X1 AOI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_10425_), .B(_10433_), .C(_10012_), .Y(_10539_) );
	XNOR2X1 XNOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_10539_), .B(_9991_), .Y(_10540_) );
	NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_9987_), .B(divider_divuResult_0_bF_buf1), .Y(_10541_) );
	AOI21X1 AOI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf0), .B(_10540_), .C(_10541_), .Y(divider_flipSign_rem_operand_18_) );
	OAI21X1 OAI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_9965_), .B(divider_divuResult_1_bF_buf0), .C(_9974_), .Y(_10542_) );
	NAND2X1 NAND2X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_9983_), .B(_9975_), .Y(_10543_) );
	OAI21X1 OAI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_9991_), .B(_10539_), .C(_9988_), .Y(_10545_) );
	OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_10545_), .B(_10543_), .Y(_10546_) );
	NAND2X1 NAND2X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_10543_), .B(_10545_), .Y(_10547_) );
	NAND3X1 NAND3X1_2233 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf6), .B(_10547_), .C(_10546_), .Y(_10548_) );
	OAI21X1 OAI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_10542_), .B(divider_divuResult_0_bF_buf5), .C(_10548_), .Y(divider_flipSign_rem_operand_19_) );
	INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(_10017_), .Y(_10549_) );
	AOI21X1 AOI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(_10424_), .C(_10434_), .Y(_10550_) );
	OAI21X1 OAI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_10549_), .B(_10550_), .C(_9961_), .Y(_10551_) );
	INVX1 INVX1_1439 ( .gnd(gnd), .vdd(vdd), .A(_9961_), .Y(_10552_) );
	AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_10433_), .B(_9993_), .Y(_10553_) );
	AOI21X1 AOI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_10425_), .B(_10553_), .C(_10549_), .Y(_10555_) );
	NAND2X1 NAND2X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_10552_), .B(_10555_), .Y(_10556_) );
	NAND3X1 NAND3X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_10551_), .B(_10556_), .C(divider_divuResult_0_bF_buf4), .Y(_10557_) );
	OAI21X1 OAI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_10018_), .B(divider_divuResult_0_bF_buf3), .C(_10557_), .Y(divider_flipSign_rem_operand_20_) );
	OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_9955_), .B(_4424__bF_buf1), .Y(_10558_) );
	NAND2X1 NAND2X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_4424__bF_buf0), .B(_9955_), .Y(_10559_) );
	NAND2X1 NAND2X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_10559_), .B(_10558_), .Y(_10560_) );
	NAND2X1 NAND2X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_4011__bF_buf3), .B(_9960_), .Y(_10561_) );
	OAI21X1 OAI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_10552_), .B(_10555_), .C(_10561_), .Y(_10562_) );
	XNOR2X1 XNOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_10562_), .B(_10560_), .Y(_10563_) );
	MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_10563_), .B(_9955_), .S(divider_divuResult_0_bF_buf2), .Y(divider_flipSign_rem_operand_21_) );
	INVX1 INVX1_1440 ( .gnd(gnd), .vdd(vdd), .A(_9938_), .Y(_10565_) );
	NAND3X1 NAND3X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_10226_), .B(_10253_), .C(_10458_), .Y(_10566_) );
	INVX1 INVX1_1441 ( .gnd(gnd), .vdd(vdd), .A(_10403_), .Y(_10567_) );
	NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_10488_), .B(_10406_), .Y(_10568_) );
	NAND3X1 NAND3X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_10567_), .B(_10336_), .C(_10568_), .Y(_10569_) );
	AOI21X1 AOI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_10566_), .B(_10260_), .C(_10569_), .Y(_10570_) );
	INVX1 INVX1_1442 ( .gnd(gnd), .vdd(vdd), .A(_10423_), .Y(_10571_) );
	OAI21X1 OAI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_10337_), .B(_10502_), .C(_10571_), .Y(_10572_) );
	OAI21X1 OAI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_10572_), .B(_10570_), .C(_10553_), .Y(_10573_) );
	AOI21X1 AOI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_10573_), .B(_10017_), .C(_9962_), .Y(_10575_) );
	OAI21X1 OAI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_10021_), .B(_10575_), .C(_10426_), .Y(_10576_) );
	INVX1 INVX1_1443 ( .gnd(gnd), .vdd(vdd), .A(_10426_), .Y(_10577_) );
	OAI21X1 OAI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_10549_), .B(_10550_), .C(_9963_), .Y(_10578_) );
	NAND3X1 NAND3X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_10577_), .B(_10020_), .C(_10578_), .Y(_10579_) );
	NAND3X1 NAND3X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_10576_), .B(_10579_), .C(divider_divuResult_0_bF_buf1), .Y(_10580_) );
	OAI21X1 OAI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_10565_), .B(divider_divuResult_0_bF_buf0), .C(_10580_), .Y(divider_flipSign_rem_operand_22_) );
	OAI21X1 OAI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_9928_), .B(divider_divuResult_1_bF_buf6), .C(_9925_), .Y(_10581_) );
	OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf6), .B(_10581_), .Y(_10582_) );
	NAND2X1 NAND2X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_9927_), .B(_9933_), .Y(_10583_) );
	INVX1 INVX1_1444 ( .gnd(gnd), .vdd(vdd), .A(_10583_), .Y(_10585_) );
	NAND3X1 NAND3X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_10585_), .B(_10024_), .C(_10576_), .Y(_10586_) );
	AOI21X1 AOI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_10578_), .B(_10020_), .C(_10577_), .Y(_10587_) );
	OAI21X1 OAI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_10026_), .B(_10587_), .C(_10583_), .Y(_10588_) );
	NAND3X1 NAND3X1_2240 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf5), .B(_10586_), .C(_10588_), .Y(_10589_) );
	NAND2X1 NAND2X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_10582_), .B(_10589_), .Y(divider_flipSign_rem_operand_23_) );
	INVX1 INVX1_1445 ( .gnd(gnd), .vdd(vdd), .A(_10145_), .Y(_10590_) );
	NAND3X1 NAND3X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_9943_), .B(_9963_), .C(_10553_), .Y(_10591_) );
	AOI21X1 AOI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(_10424_), .C(_10591_), .Y(_10592_) );
	OAI21X1 OAI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_10030_), .B(_10592_), .C(_10590_), .Y(_10593_) );
	NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_9962_), .B(_10427_), .Y(_10595_) );
	INVX1 INVX1_1446 ( .gnd(gnd), .vdd(vdd), .A(_10022_), .Y(_10596_) );
	AOI21X1 AOI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_10026_), .B(_10023_), .C(_10596_), .Y(_10597_) );
	OAI21X1 OAI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_10020_), .B(_10427_), .C(_10597_), .Y(_10598_) );
	AOI21X1 AOI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_10549_), .B(_10595_), .C(_10598_), .Y(_10599_) );
	OAI21X1 OAI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_10572_), .B(_10570_), .C(_10435_), .Y(_10600_) );
	NAND3X1 NAND3X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_10145_), .B(_10599_), .C(_10600_), .Y(_10601_) );
	NAND3X1 NAND3X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_10593_), .B(_10601_), .C(divider_divuResult_0_bF_buf4), .Y(_10602_) );
	OAI21X1 OAI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_10143_), .B(divider_divuResult_0_bF_buf3), .C(_10602_), .Y(divider_flipSign_rem_operand_24_) );
	OAI21X1 OAI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_24_bF_buf3), .B(_10143_), .C(_10593_), .Y(_10603_) );
	AOI21X1 AOI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_10140_), .B(_10142_), .C(_10603_), .Y(_10605_) );
	INVX1 INVX1_1447 ( .gnd(gnd), .vdd(vdd), .A(_10072_), .Y(_10606_) );
	AOI22X1 AOI22X1_234 ( .gnd(gnd), .vdd(vdd), .A(_10606_), .B(_10073_), .C(_10079_), .D(_10593_), .Y(_10607_) );
	OAI21X1 OAI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_10607_), .B(_10605_), .C(divider_divuResult_0_bF_buf2), .Y(_10608_) );
	OAI21X1 OAI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_10141_), .B(divider_divuResult_0_bF_buf1), .C(_10608_), .Y(divider_flipSign_rem_operand_25_) );
	NAND2X1 NAND2X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_10056_), .B(_10057_), .Y(_10609_) );
	INVX1 INVX1_1448 ( .gnd(gnd), .vdd(vdd), .A(_10147_), .Y(_10610_) );
	AOI21X1 AOI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_10600_), .B(_10599_), .C(_10610_), .Y(_10611_) );
	OAI21X1 OAI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_10081_), .B(_10611_), .C(_10609_), .Y(_10612_) );
	INVX1 INVX1_1449 ( .gnd(gnd), .vdd(vdd), .A(_10609_), .Y(_10613_) );
	INVX1 INVX1_1450 ( .gnd(gnd), .vdd(vdd), .A(_10081_), .Y(_10614_) );
	OAI21X1 OAI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_10030_), .B(_10592_), .C(_10147_), .Y(_10615_) );
	NAND3X1 NAND3X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_10613_), .B(_10614_), .C(_10615_), .Y(_10616_) );
	NAND2X1 NAND2X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_10616_), .B(_10612_), .Y(_10617_) );
	NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_10055_), .B(divider_divuResult_0_bF_buf0), .Y(_10618_) );
	AOI21X1 AOI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf6), .B(_10617_), .C(_10618_), .Y(divider_flipSign_rem_operand_26_) );
	OAI21X1 OAI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_10045_), .B(divider_divuResult_1_bF_buf5), .C(_10043_), .Y(_10619_) );
	OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf5), .B(_10619_), .Y(_10620_) );
	NAND2X1 NAND2X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_10044_), .B(_10051_), .Y(_10621_) );
	INVX1 INVX1_1451 ( .gnd(gnd), .vdd(vdd), .A(_10621_), .Y(_10622_) );
	NAND3X1 NAND3X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_10622_), .B(_10084_), .C(_10612_), .Y(_10624_) );
	INVX1 INVX1_1452 ( .gnd(gnd), .vdd(vdd), .A(_10084_), .Y(_10625_) );
	AOI21X1 AOI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_10615_), .B(_10614_), .C(_10613_), .Y(_10626_) );
	OAI21X1 OAI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_10625_), .B(_10626_), .C(_10621_), .Y(_10627_) );
	NAND3X1 NAND3X1_2246 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf4), .B(_10624_), .C(_10627_), .Y(_10628_) );
	NAND2X1 NAND2X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_10620_), .B(_10628_), .Y(divider_flipSign_rem_operand_27_) );
	INVX1 INVX1_1453 ( .gnd(gnd), .vdd(vdd), .A(_10086_), .Y(_10629_) );
	AOI21X1 AOI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_10600_), .B(_10599_), .C(_10148_), .Y(_10630_) );
	OAI21X1 OAI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_10629_), .B(_10630_), .C(_10115_), .Y(_10631_) );
	INVX1 INVX1_1454 ( .gnd(gnd), .vdd(vdd), .A(_10115_), .Y(_10632_) );
	INVX1 INVX1_1455 ( .gnd(gnd), .vdd(vdd), .A(_10148_), .Y(_10634_) );
	OAI21X1 OAI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_10030_), .B(_10592_), .C(_10634_), .Y(_10635_) );
	NAND3X1 NAND3X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_10632_), .B(_10086_), .C(_10635_), .Y(_10636_) );
	NAND3X1 NAND3X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10636_), .C(divider_divuResult_0_bF_buf3), .Y(_10637_) );
	OAI21X1 OAI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_10112_), .B(divider_divuResult_0_bF_buf2), .C(_10637_), .Y(divider_flipSign_rem_operand_28_) );
	OAI21X1 OAI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_10087_), .B(divider_divuResult_1_bF_buf4), .C(_10097_), .Y(_10638_) );
	OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf1), .B(_10638_), .Y(_10639_) );
	INVX1 INVX1_1456 ( .gnd(gnd), .vdd(vdd), .A(_10105_), .Y(_10640_) );
	NAND3X1 NAND3X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10640_), .C(_10631_), .Y(_10641_) );
	INVX1 INVX1_1457 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .Y(_10642_) );
	AOI21X1 AOI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_10635_), .B(_10086_), .C(_10632_), .Y(_10644_) );
	OAI21X1 OAI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_10642_), .B(_10644_), .C(_10105_), .Y(_10645_) );
	NAND3X1 NAND3X1_2250 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf0), .B(_10641_), .C(_10645_), .Y(_10646_) );
	NAND2X1 NAND2X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_10639_), .B(_10646_), .Y(divider_flipSign_rem_operand_29_) );
	NAND2X1 NAND2X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_10128_), .B(_10129_), .Y(_10647_) );
	NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_10632_), .B(_10640_), .Y(_10648_) );
	INVX1 INVX1_1458 ( .gnd(gnd), .vdd(vdd), .A(_10648_), .Y(_10649_) );
	AOI21X1 AOI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_10635_), .B(_10086_), .C(_10649_), .Y(_10650_) );
	OAI21X1 OAI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_10137_), .B(_10650_), .C(_10647_), .Y(_10651_) );
	INVX1 INVX1_1459 ( .gnd(gnd), .vdd(vdd), .A(_10647_), .Y(_10652_) );
	INVX1 INVX1_1460 ( .gnd(gnd), .vdd(vdd), .A(_10137_), .Y(_10654_) );
	OAI21X1 OAI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_10629_), .B(_10630_), .C(_10648_), .Y(_10655_) );
	NAND3X1 NAND3X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_10652_), .B(_10654_), .C(_10655_), .Y(_10656_) );
	NAND3X1 NAND3X1_2252 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf6), .B(_10656_), .C(_10651_), .Y(_10657_) );
	NAND3X1 NAND3X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_10127_), .B(_10436_), .C(_10150_), .Y(_10658_) );
	NAND2X1 NAND2X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_10658_), .B(_10657_), .Y(divider_flipSign_rem_operand_30_) );
	NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_1878_), .B(_2283_), .Y(_10659_) );
	XNOR2X1 XNOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_10659_), .B(_1867_), .Y(_10660_) );
	NAND2X1 NAND2X1_1815 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_30_), .B(_10660_), .Y(_10661_) );
	OAI21X1 OAI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_10118_), .B(divider_divuResult_0_bF_buf5), .C(_10661_), .Y(divider_flipSign_rem_operand_31_) );
	XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(divider_a_isNegative_bF_buf8), .Y(divider_divFlip) );
	AOI21X1 AOI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_result_0_bF_buf1), .B(_2251_), .C(_1823_), .Y(divider_divuResult_31_) );
	INVX1 INVX1_1461 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .Y(_10684_) );
	NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(comparator_unsignedEn), .B(_10684_), .Y(divider_a_isNegative) );
	INVX8 INVX8_41 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf7), .Y(_10855_) );
	NAND2X1 NAND2X1_1816 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf4), .B(_10855__bF_buf4), .Y(_10856_) );
	XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(aOperand_frameOut_0_bF_buf3), .Y(_10857_) );
	XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(aOperand_frameOut_1_bF_buf3), .Y(_10858_) );
	NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_10857_), .B(_10858_), .Y(_10859_) );
	OAI21X1 OAI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf2), .B(aOperand_frameOut_1_bF_buf2), .C(divider_a_isNegative_bF_buf4), .Y(_10860_) );
	OAI21X1 OAI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_10860_), .B(_10859_), .C(_10856_), .Y(divider_aOp_abs_1_) );
	INVX1 INVX1_1462 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf3), .Y(_10861_) );
	AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_10857_), .B(_10858_), .Y(_10862_) );
	INVX1 INVX1_1463 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .Y(_10863_) );
	OAI21X1 OAI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf2), .B(_10863_), .C(divider_a_isNegative_bF_buf3), .Y(_10864_) );
	NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_10861_), .B(_10862_), .Y(_10865_) );
	OAI22X1 OAI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(_10861_), .C(_10865_), .D(_10864_), .Y(divider_aOp_abs_2_) );
	XNOR2X1 XNOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_10864_), .B(aOperand_frameOut_3_bF_buf4), .Y(divider_aOp_abs_3_) );
	NAND2X1 NAND2X1_1817 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf4), .B(_10855__bF_buf3), .Y(_10866_) );
	NAND3X1 NAND3X1_2254 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf1), .B(aOperand_frameOut_3_bF_buf3), .C(_10855__bF_buf2), .Y(_10867_) );
	INVX1 INVX1_1464 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .Y(_10868_) );
	NAND3X1 NAND3X1_2255 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(_10861_), .C(_10868_), .Y(_10869_) );
	NAND2X1 NAND2X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_10867_), .B(_10869_), .Y(_10870_) );
	NAND3X1 NAND3X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_10857_), .B(_10858_), .C(_10870_), .Y(_10871_) );
	INVX1 INVX1_1465 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .Y(_10872_) );
	NAND2X1 NAND2X1_1819 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(_10872_), .Y(_10873_) );
	NAND2X1 NAND2X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_10866_), .B(_10873_), .Y(_10874_) );
	XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_10871_), .B(_10874_), .Y(_10875_) );
	OAI21X1 OAI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_10855__bF_buf1), .B(_10875_), .C(_10866_), .Y(divider_aOp_abs_4_) );
	INVX1 INVX1_1466 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf3), .Y(_10876_) );
	NAND3X1 NAND3X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_10870_), .B(_10874_), .C(_10862_), .Y(_10877_) );
	NAND2X1 NAND2X1_1821 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf2), .B(_10855__bF_buf0), .Y(_10878_) );
	NAND2X1 NAND2X1_1822 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf8), .B(_10876_), .Y(_10879_) );
	NAND2X1 NAND2X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_10878_), .B(_10879_), .Y(_10880_) );
	NAND2X1 NAND2X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .B(_10877_), .Y(_10881_) );
	OAI21X1 OAI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_10876_), .B(_10877_), .C(_10881_), .Y(divider_aOp_abs_5_) );
	OAI21X1 OAI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf1), .B(_10877_), .C(divider_a_isNegative_bF_buf7), .Y(_10882_) );
	XNOR2X1 XNOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_10882_), .B(aOperand_frameOut_6_bF_buf0), .Y(divider_aOp_abs_6_) );
	INVX1 INVX1_1467 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf4), .Y(_10685_) );
	AOI21X1 AOI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_10878_), .B(_10879_), .C(_10877_), .Y(_10686_) );
	NAND2X1 NAND2X1_1825 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf4), .B(_10855__bF_buf4), .Y(_10687_) );
	INVX1 INVX1_1468 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf3), .Y(_10688_) );
	NAND2X1 NAND2X1_1826 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(_10688_), .Y(_10689_) );
	NAND2X1 NAND2X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_10687_), .B(_10689_), .Y(_10690_) );
	NAND2X1 NAND2X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_10690_), .B(_10686_), .Y(_10691_) );
	NAND2X1 NAND2X1_1829 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf3), .B(_10855__bF_buf3), .Y(_10692_) );
	NAND2X1 NAND2X1_1830 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(_10685_), .Y(_10693_) );
	NAND2X1 NAND2X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_10692_), .B(_10693_), .Y(_10694_) );
	NAND2X1 NAND2X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_10694_), .B(_10691_), .Y(_10695_) );
	OAI21X1 OAI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_10685_), .B(_10691_), .C(_10695_), .Y(divider_aOp_abs_7_) );
	AOI22X1 AOI22X1_235 ( .gnd(gnd), .vdd(vdd), .A(_10866_), .B(_10873_), .C(_10878_), .D(_10879_), .Y(_10696_) );
	AOI22X1 AOI22X1_236 ( .gnd(gnd), .vdd(vdd), .A(_10687_), .B(_10689_), .C(_10692_), .D(_10693_), .Y(_10697_) );
	NAND2X1 NAND2X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_10696_), .B(_10697_), .Y(_10698_) );
	OAI21X1 OAI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_10871_), .B(_10698_), .C(divider_a_isNegative_bF_buf4), .Y(_10699_) );
	XNOR2X1 XNOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_10699_), .B(aOperand_frameOut_8_bF_buf4), .Y(divider_aOp_abs_8_) );
	INVX1 INVX1_1469 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf3), .Y(_10700_) );
	NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_10871_), .B(_10698_), .Y(_10701_) );
	NAND2X1 NAND2X1_1834 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf3), .B(_10855__bF_buf2), .Y(_10702_) );
	INVX1 INVX1_1470 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf2), .Y(_10703_) );
	NAND2X1 NAND2X1_1835 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(_10703_), .Y(_10704_) );
	NAND2X1 NAND2X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_10702_), .B(_10704_), .Y(_10705_) );
	NAND2X1 NAND2X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_10705_), .B(_10701_), .Y(_10706_) );
	NAND2X1 NAND2X1_1838 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf2), .B(_10855__bF_buf1), .Y(_10707_) );
	NAND2X1 NAND2X1_1839 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(_10700_), .Y(_10708_) );
	NAND2X1 NAND2X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_10707_), .B(_10708_), .Y(_10709_) );
	NAND2X1 NAND2X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_10709_), .B(_10706_), .Y(_10710_) );
	OAI21X1 OAI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_10700_), .B(_10706_), .C(_10710_), .Y(divider_aOp_abs_9_) );
	OAI21X1 OAI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf1), .B(_10706_), .C(divider_a_isNegative_bF_buf1), .Y(_10711_) );
	XNOR2X1 XNOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_10711_), .B(aOperand_frameOut_10_bF_buf4), .Y(divider_aOp_abs_10_) );
	INVX1 INVX1_1471 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf0), .Y(_10712_) );
	AOI22X1 AOI22X1_237 ( .gnd(gnd), .vdd(vdd), .A(_10702_), .B(_10704_), .C(_10707_), .D(_10708_), .Y(_10713_) );
	NAND2X1 NAND2X1_1842 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf3), .B(_10855__bF_buf0), .Y(_10714_) );
	INVX1 INVX1_1472 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf2), .Y(_10715_) );
	NAND2X1 NAND2X1_1843 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(_10715_), .Y(_10716_) );
	NAND2X1 NAND2X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_10714_), .B(_10716_), .Y(_10717_) );
	NAND3X1 NAND3X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_10713_), .B(_10717_), .C(_10701_), .Y(_10718_) );
	NAND2X1 NAND2X1_1845 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf4), .B(_10855__bF_buf4), .Y(_10719_) );
	NAND2X1 NAND2X1_1846 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf8), .B(_10712_), .Y(_10720_) );
	NAND2X1 NAND2X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_10719_), .B(_10720_), .Y(_10721_) );
	NAND2X1 NAND2X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_10721_), .B(_10718_), .Y(_10722_) );
	OAI21X1 OAI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_10712_), .B(_10718_), .C(_10722_), .Y(divider_aOp_abs_11_) );
	NAND2X1 NAND2X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_10713_), .B(_10701_), .Y(_10723_) );
	AOI22X1 AOI22X1_238 ( .gnd(gnd), .vdd(vdd), .A(_10714_), .B(_10716_), .C(_10719_), .D(_10720_), .Y(_10724_) );
	INVX1 INVX1_1473 ( .gnd(gnd), .vdd(vdd), .A(_10724_), .Y(_10725_) );
	OAI21X1 OAI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_10725_), .B(_10723_), .C(divider_a_isNegative_bF_buf7), .Y(_10726_) );
	XNOR2X1 XNOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_10726_), .B(aOperand_frameOut_12_bF_buf4), .Y(divider_aOp_abs_12_) );
	INVX1 INVX1_1474 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf3), .Y(_10727_) );
	NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_10725_), .B(_10723_), .Y(_10728_) );
	NAND2X1 NAND2X1_1850 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf3), .B(_10855__bF_buf3), .Y(_10729_) );
	INVX1 INVX1_1475 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf2), .Y(_10730_) );
	NAND2X1 NAND2X1_1851 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(_10730_), .Y(_10731_) );
	NAND2X1 NAND2X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_10729_), .B(_10731_), .Y(_10732_) );
	NAND2X1 NAND2X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_10732_), .B(_10728_), .Y(_10733_) );
	NAND2X1 NAND2X1_1854 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf2), .B(_10855__bF_buf2), .Y(_10734_) );
	NAND2X1 NAND2X1_1855 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(_10727_), .Y(_10735_) );
	NAND2X1 NAND2X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_10734_), .B(_10735_), .Y(_10736_) );
	NAND2X1 NAND2X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_10736_), .B(_10733_), .Y(_10737_) );
	OAI21X1 OAI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_10727_), .B(_10733_), .C(_10737_), .Y(divider_aOp_abs_13_) );
	INVX1 INVX1_1476 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf4), .Y(_10738_) );
	NAND3X1 NAND3X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_10713_), .B(_10724_), .C(_10701_), .Y(_10739_) );
	AOI22X1 AOI22X1_239 ( .gnd(gnd), .vdd(vdd), .A(_10729_), .B(_10731_), .C(_10734_), .D(_10735_), .Y(_10740_) );
	INVX1 INVX1_1477 ( .gnd(gnd), .vdd(vdd), .A(_10740_), .Y(_10741_) );
	NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_10741_), .B(_10739_), .Y(_10742_) );
	NAND2X1 NAND2X1_1858 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf3), .B(_10855__bF_buf1), .Y(_10743_) );
	NAND2X1 NAND2X1_1859 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(_10738_), .Y(_10744_) );
	NAND2X1 NAND2X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_10743_), .B(_10744_), .Y(_10745_) );
	AOI21X1 AOI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_10728_), .B(_10740_), .C(_10745_), .Y(_10746_) );
	AOI21X1 AOI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_10738_), .B(_10742_), .C(_10746_), .Y(divider_aOp_abs_14_) );
	INVX1 INVX1_1478 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf4), .Y(_10747_) );
	NAND2X1 NAND2X1_1861 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf3), .B(_10855__bF_buf0), .Y(_10748_) );
	NAND2X1 NAND2X1_1862 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(_10747_), .Y(_10749_) );
	NAND2X1 NAND2X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_10748_), .B(_10749_), .Y(_10750_) );
	INVX1 INVX1_1479 ( .gnd(gnd), .vdd(vdd), .A(_10750_), .Y(_10751_) );
	NAND2X1 NAND2X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_10745_), .B(_10742_), .Y(_10752_) );
	MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_10751_), .B(_10747_), .S(_10752_), .Y(divider_aOp_abs_15_) );
	NAND2X1 NAND2X1_1865 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf3), .B(_10855__bF_buf4), .Y(_10753_) );
	NAND2X1 NAND2X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_10713_), .B(_10724_), .Y(_10754_) );
	AOI22X1 AOI22X1_240 ( .gnd(gnd), .vdd(vdd), .A(_10743_), .B(_10744_), .C(_10748_), .D(_10749_), .Y(_10755_) );
	NAND2X1 NAND2X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_10740_), .B(_10755_), .Y(_10756_) );
	NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_10754_), .B(_10756_), .Y(_10757_) );
	AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_10757_), .B(_10701_), .Y(_10758_) );
	INVX1 INVX1_1480 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf2), .Y(_10759_) );
	NAND2X1 NAND2X1_1868 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(_10759_), .Y(_10760_) );
	NAND2X1 NAND2X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_10753_), .B(_10760_), .Y(_10761_) );
	XNOR2X1 XNOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_10758_), .B(_10761_), .Y(_10762_) );
	OAI21X1 OAI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_10855__bF_buf3), .B(_10762_), .C(_10753_), .Y(divider_aOp_abs_16_) );
	INVX1 INVX1_1481 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf4), .Y(_10763_) );
	NAND2X1 NAND2X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_10713_), .B(_10755_), .Y(_10764_) );
	NAND2X1 NAND2X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_10724_), .B(_10740_), .Y(_10765_) );
	NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_10764_), .B(_10765_), .Y(_10766_) );
	AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_10766_), .B(_10701_), .Y(_10767_) );
	NAND2X1 NAND2X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_10761_), .B(_10767_), .Y(_10768_) );
	INVX1 INVX1_1482 ( .gnd(gnd), .vdd(vdd), .A(_10758_), .Y(_10769_) );
	INVX1 INVX1_1483 ( .gnd(gnd), .vdd(vdd), .A(_10761_), .Y(_10770_) );
	NAND2X1 NAND2X1_1873 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf3), .B(_10855__bF_buf2), .Y(_10771_) );
	NAND2X1 NAND2X1_1874 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(_10763_), .Y(_10772_) );
	NAND2X1 NAND2X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_10771_), .B(_10772_), .Y(_10773_) );
	OAI21X1 OAI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_10770_), .B(_10769_), .C(_10773_), .Y(_10774_) );
	OAI21X1 OAI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_10763_), .B(_10768_), .C(_10774_), .Y(divider_aOp_abs_17_) );
	INVX1 INVX1_1484 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf3), .Y(_10775_) );
	AOI22X1 AOI22X1_241 ( .gnd(gnd), .vdd(vdd), .A(_10753_), .B(_10760_), .C(_10771_), .D(_10772_), .Y(_10776_) );
	AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_10767_), .B(_10776_), .Y(_10777_) );
	NAND2X1 NAND2X1_1876 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf2), .B(_10855__bF_buf1), .Y(_10778_) );
	NAND2X1 NAND2X1_1877 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(_10775_), .Y(_10779_) );
	NAND2X1 NAND2X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_10778_), .B(_10779_), .Y(_10780_) );
	NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_10780_), .B(_10777_), .Y(_10781_) );
	AOI21X1 AOI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_10775_), .B(_10777_), .C(_10781_), .Y(divider_aOp_abs_18_) );
	INVX1 INVX1_1485 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf3), .Y(_10782_) );
	NAND2X1 NAND2X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_10780_), .B(_10777_), .Y(_10783_) );
	XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf8), .B(aOperand_frameOut_19_bF_buf2), .Y(_10784_) );
	NAND2X1 NAND2X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_10784_), .B(_10783_), .Y(_10785_) );
	OAI21X1 OAI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_10782_), .B(_10783_), .C(_10785_), .Y(divider_aOp_abs_19_) );
	NAND3X1 NAND3X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_10780_), .B(_10784_), .C(_10776_), .Y(_10786_) );
	OAI21X1 OAI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10769_), .C(divider_a_isNegative_bF_buf7), .Y(_10787_) );
	XNOR2X1 XNOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_10787_), .B(aOperand_frameOut_20_bF_buf0), .Y(divider_aOp_abs_20_) );
	INVX1 INVX1_1486 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf2), .Y(_10788_) );
	NAND2X1 NAND2X1_1881 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf1), .B(_10855__bF_buf0), .Y(_10789_) );
	NAND2X1 NAND2X1_1882 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(_10788_), .Y(_10790_) );
	AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_10789_), .B(_10790_), .Y(_10791_) );
	INVX1 INVX1_1487 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .Y(_10792_) );
	NAND2X1 NAND2X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_10792_), .B(_10767_), .Y(_10793_) );
	NAND2X1 NAND2X1_1884 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf4), .B(_10855__bF_buf4), .Y(_10794_) );
	INVX1 INVX1_1488 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf3), .Y(_10795_) );
	NAND2X1 NAND2X1_1885 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(_10795_), .Y(_10796_) );
	AOI21X1 AOI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_10794_), .B(_10796_), .C(_10793_), .Y(_10797_) );
	MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_10788_), .B(_10791_), .S(_10797_), .Y(divider_aOp_abs_21_) );
	INVX1 INVX1_1489 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf3), .Y(_10798_) );
	NAND2X1 NAND2X1_1886 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf2), .B(_10855__bF_buf3), .Y(_10799_) );
	NAND2X1 NAND2X1_1887 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(_10798_), .Y(_10800_) );
	NAND2X1 NAND2X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_10799_), .B(_10800_), .Y(_10801_) );
	INVX1 INVX1_1490 ( .gnd(gnd), .vdd(vdd), .A(_10801_), .Y(_10802_) );
	AOI22X1 AOI22X1_242 ( .gnd(gnd), .vdd(vdd), .A(_10794_), .B(_10796_), .C(_10789_), .D(_10790_), .Y(_10803_) );
	INVX1 INVX1_1491 ( .gnd(gnd), .vdd(vdd), .A(_10803_), .Y(_10804_) );
	NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_10804_), .B(_10793_), .Y(_10805_) );
	MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .B(_10802_), .S(_10805_), .Y(divider_aOp_abs_22_) );
	XOR2X1 XOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(aOperand_frameOut_23_), .Y(_10806_) );
	INVX1 INVX1_1492 ( .gnd(gnd), .vdd(vdd), .A(_10806_), .Y(_10807_) );
	NAND2X1 NAND2X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_10792_), .B(_10758_), .Y(_10808_) );
	NOR3X1 NOR3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_10802_), .B(_10804_), .C(_10808_), .Y(_10809_) );
	NAND3X1 NAND3X1_2261 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .B(_10801_), .C(_10805_), .Y(_10810_) );
	OAI21X1 OAI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_10807_), .B(_10809_), .C(_10810_), .Y(divider_aOp_abs_23_) );
	NAND2X1 NAND2X1_1890 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf2), .B(_10855__bF_buf2), .Y(_10811_) );
	INVX1 INVX1_1493 ( .gnd(gnd), .vdd(vdd), .A(_10811_), .Y(_10812_) );
	NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf1), .B(_10855__bF_buf1), .Y(_10813_) );
	OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_10812_), .B(_10813_), .Y(_10814_) );
	NAND3X1 NAND3X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_10801_), .B(_10806_), .C(_10803_), .Y(_10815_) );
	NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_10786_), .B(_10815_), .Y(_10816_) );
	NAND3X1 NAND3X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_10701_), .B(_10757_), .C(_10816_), .Y(_10817_) );
	XOR2X1 XOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_10817_), .B(_10814_), .Y(_10818_) );
	OAI21X1 OAI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_10855__bF_buf0), .B(_10818_), .C(_10811_), .Y(divider_aOp_abs_24_) );
	OAI21X1 OAI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf0), .B(_10817_), .C(divider_a_isNegative_bF_buf2), .Y(_10819_) );
	XNOR2X1 XNOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_10819_), .B(aOperand_frameOut_25_bF_buf2), .Y(divider_aOp_abs_25_) );
	XOR2X1 XOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(aOperand_frameOut_25_bF_buf1), .Y(_10820_) );
	OAI21X1 OAI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_10813_), .B(_10812_), .C(_10820_), .Y(_10821_) );
	OAI21X1 OAI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .B(_10817_), .C(divider_a_isNegative_bF_buf0), .Y(_10822_) );
	XNOR2X1 XNOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_10822_), .B(aOperand_frameOut_26_), .Y(divider_aOp_abs_26_) );
	XOR2X1 XOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf8), .B(aOperand_frameOut_27_), .Y(_10823_) );
	INVX1 INVX1_1494 ( .gnd(gnd), .vdd(vdd), .A(_10823_), .Y(_10824_) );
	NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .B(_10817_), .Y(_10825_) );
	XOR2X1 XOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf7), .B(aOperand_frameOut_26_), .Y(_10826_) );
	NAND2X1 NAND2X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_10826_), .B(_10825_), .Y(_10827_) );
	NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_27_), .B(_10827_), .Y(_10828_) );
	AOI21X1 AOI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_10824_), .B(_10827_), .C(_10828_), .Y(divider_aOp_abs_27_) );
	INVX1 INVX1_1495 ( .gnd(gnd), .vdd(vdd), .A(_10821_), .Y(_10829_) );
	AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_10826_), .B(_10823_), .Y(_10830_) );
	NAND2X1 NAND2X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_10830_), .B(_10829_), .Y(_10831_) );
	OAI21X1 OAI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .B(_10817_), .C(divider_a_isNegative_bF_buf6), .Y(_10832_) );
	XNOR2X1 XNOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_10832_), .B(aOperand_frameOut_28_), .Y(divider_aOp_abs_28_) );
	XOR2X1 XOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(aOperand_frameOut_29_), .Y(_10833_) );
	INVX1 INVX1_1496 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .Y(_10834_) );
	NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .B(_10817_), .Y(_10835_) );
	XNOR2X1 XNOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(aOperand_frameOut_28_), .Y(_10836_) );
	INVX1 INVX1_1497 ( .gnd(gnd), .vdd(vdd), .A(_10836_), .Y(_10837_) );
	NAND2X1 NAND2X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_10837_), .B(_10835_), .Y(_10838_) );
	NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .B(_10838_), .Y(_10839_) );
	AOI21X1 AOI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_10834_), .B(_10838_), .C(_10839_), .Y(divider_aOp_abs_29_) );
	INVX1 INVX1_1498 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .Y(_10840_) );
	NAND2X1 NAND2X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .B(_10837_), .Y(_10841_) );
	NOR3X1 NOR3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .B(_10841_), .C(_10817_), .Y(_10842_) );
	OAI21X1 OAI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_10855__bF_buf4), .B(_10842_), .C(_10840_), .Y(_10843_) );
	INVX1 INVX1_1499 ( .gnd(gnd), .vdd(vdd), .A(_10841_), .Y(_10844_) );
	NAND2X1 NAND2X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_10844_), .B(_10835_), .Y(_10845_) );
	NAND3X1 NAND3X1_2264 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(aOperand_frameOut_30_), .C(_10845_), .Y(_10846_) );
	AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_10846_), .B(_10843_), .Y(divider_aOp_abs_30_) );
	INVX1 INVX1_1500 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .Y(_10847_) );
	NAND3X1 NAND3X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_10840_), .B(_10844_), .C(_10835_), .Y(_10848_) );
	NAND3X1 NAND3X1_2266 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(_10847_), .C(_10848_), .Y(_10849_) );
	INVX1 INVX1_1501 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .Y(_10850_) );
	NAND3X1 NAND3X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_10816_), .B(_10850_), .C(_10758_), .Y(_10851_) );
	OAI21X1 OAI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_10841_), .B(_10851_), .C(divider_a_isNegative_bF_buf1), .Y(_10852_) );
	NAND2X1 NAND2X1_1896 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(aOperand_frameOut_30_), .Y(_10853_) );
	NAND3X1 NAND3X1_2268 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .B(_10853_), .C(_10852_), .Y(_10854_) );
	NAND2X1 NAND2X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_10849_), .B(_10854_), .Y(divider_aOp_abs_31_) );
	BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf1), .Y(divider_aOp_abs_0_) );
	INVX1 INVX1_1502 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_msb), .Y(_10883_) );
	NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(comparator_unsignedEn), .B(_10883_), .Y(divider_absoluteValue_B_flipSign_flip) );
	INVX8 INVX8_42 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf4), .Y(_11054_) );
	NAND2X1 NAND2X1_1898 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf1), .B(_11054__bF_buf4), .Y(_11055_) );
	XOR2X1 XOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(adder_bOperand_0_bF_buf2), .Y(_11056_) );
	XOR2X1 XOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf2), .B(adder_bOperand_1_bF_buf0), .Y(_11057_) );
	NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_11056_), .B(_11057_), .Y(_11058_) );
	OAI21X1 OAI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(adder_bOperand_1_bF_buf6), .C(divider_absoluteValue_B_flipSign_flip_bF_buf1), .Y(_11059_) );
	OAI21X1 OAI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_11059_), .B(_11058_), .C(_11055_), .Y(divider_absoluteValue_B_flipSign_result_1_) );
	INVX1 INVX1_1503 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .Y(_11060_) );
	AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_11056_), .B(_11057_), .Y(_11061_) );
	INVX1 INVX1_1504 ( .gnd(gnd), .vdd(vdd), .A(_11061_), .Y(_11062_) );
	OAI21X1 OAI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf3), .B(_11062_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf0), .Y(_11063_) );
	NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11061_), .Y(_11064_) );
	OAI22X1 OAI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(_11060_), .C(_11064_), .D(_11063_), .Y(divider_absoluteValue_B_flipSign_result_2_) );
	XNOR2X1 XNOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_11063_), .B(adder_bOperand_3_bF_buf0), .Y(divider_absoluteValue_B_flipSign_result_3_) );
	NAND2X1 NAND2X1_1899 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf0), .B(_11054__bF_buf3), .Y(_11065_) );
	NAND3X1 NAND3X1_2269 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf2), .B(adder_bOperand_3_bF_buf5), .C(_11054__bF_buf2), .Y(_11066_) );
	INVX1 INVX1_1505 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .Y(_11067_) );
	NAND3X1 NAND3X1_2270 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf4), .B(_11060_), .C(_11067_), .Y(_11068_) );
	NAND2X1 NAND2X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_11066_), .B(_11068_), .Y(_11069_) );
	NAND3X1 NAND3X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_11056_), .B(_11057_), .C(_11069_), .Y(_11070_) );
	INVX1 INVX1_1506 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf5), .Y(_11071_) );
	NAND2X1 NAND2X1_1901 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(_11071_), .Y(_11072_) );
	NAND2X1 NAND2X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_11065_), .B(_11072_), .Y(_11073_) );
	XOR2X1 XOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_11070_), .B(_11073_), .Y(_11074_) );
	OAI21X1 OAI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_11054__bF_buf1), .B(_11074_), .C(_11065_), .Y(divider_absoluteValue_B_flipSign_result_4_) );
	INVX1 INVX1_1507 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf4), .Y(_11075_) );
	NAND3X1 NAND3X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .B(_11073_), .C(_11061_), .Y(_11076_) );
	NAND2X1 NAND2X1_1903 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf3), .B(_11054__bF_buf0), .Y(_11077_) );
	NAND2X1 NAND2X1_1904 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf2), .B(_11075_), .Y(_11078_) );
	NAND2X1 NAND2X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_11077_), .B(_11078_), .Y(_11079_) );
	NAND2X1 NAND2X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_11079_), .B(_11076_), .Y(_11080_) );
	OAI21X1 OAI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_11075_), .B(_11076_), .C(_11080_), .Y(divider_absoluteValue_B_flipSign_result_5_) );
	OAI21X1 OAI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf2), .B(_11076_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf1), .Y(_11081_) );
	XNOR2X1 XNOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_11081_), .B(adder_bOperand_6_bF_buf0), .Y(divider_absoluteValue_B_flipSign_result_6_) );
	INVX1 INVX1_1508 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf0), .Y(_10884_) );
	AOI21X1 AOI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_11077_), .B(_11078_), .C(_11076_), .Y(_10885_) );
	NAND2X1 NAND2X1_1907 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(_11054__bF_buf4), .Y(_10886_) );
	INVX1 INVX1_1509 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf4), .Y(_10887_) );
	NAND2X1 NAND2X1_1908 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf0), .B(_10887_), .Y(_10888_) );
	NAND2X1 NAND2X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_10886_), .B(_10888_), .Y(_10889_) );
	NAND2X1 NAND2X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_10889_), .B(_10885_), .Y(_10890_) );
	NAND2X1 NAND2X1_1911 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(_11054__bF_buf3), .Y(_10891_) );
	NAND2X1 NAND2X1_1912 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(_10884_), .Y(_10892_) );
	NAND2X1 NAND2X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_10891_), .B(_10892_), .Y(_10893_) );
	NAND2X1 NAND2X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_10893_), .B(_10890_), .Y(_10894_) );
	OAI21X1 OAI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_10884_), .B(_10890_), .C(_10894_), .Y(divider_absoluteValue_B_flipSign_result_7_) );
	AOI22X1 AOI22X1_243 ( .gnd(gnd), .vdd(vdd), .A(_11065_), .B(_11072_), .C(_11077_), .D(_11078_), .Y(_10895_) );
	AOI22X1 AOI22X1_244 ( .gnd(gnd), .vdd(vdd), .A(_10886_), .B(_10888_), .C(_10891_), .D(_10892_), .Y(_10896_) );
	NAND2X1 NAND2X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_10895_), .B(_10896_), .Y(_10897_) );
	OAI21X1 OAI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_11070_), .B(_10897_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf4), .Y(_10898_) );
	XNOR2X1 XNOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_10898_), .B(adder_bOperand_8_bF_buf4), .Y(divider_absoluteValue_B_flipSign_result_8_) );
	INVX1 INVX1_1510 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf0), .Y(_10899_) );
	NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_11070_), .B(_10897_), .Y(_10900_) );
	NAND2X1 NAND2X1_1916 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf3), .B(_11054__bF_buf2), .Y(_10901_) );
	INVX1 INVX1_1511 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf2), .Y(_10902_) );
	NAND2X1 NAND2X1_1917 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(_10902_), .Y(_10903_) );
	NAND2X1 NAND2X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_10901_), .B(_10903_), .Y(_10904_) );
	NAND2X1 NAND2X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_10904_), .B(_10900_), .Y(_10905_) );
	NAND2X1 NAND2X1_1920 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf4), .B(_11054__bF_buf1), .Y(_10906_) );
	NAND2X1 NAND2X1_1921 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf2), .B(_10899_), .Y(_10907_) );
	NAND2X1 NAND2X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_10906_), .B(_10907_), .Y(_10908_) );
	NAND2X1 NAND2X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_10908_), .B(_10905_), .Y(_10909_) );
	OAI21X1 OAI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_10899_), .B(_10905_), .C(_10909_), .Y(divider_absoluteValue_B_flipSign_result_9_) );
	OAI21X1 OAI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf3), .B(_10905_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf1), .Y(_10910_) );
	XNOR2X1 XNOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_10910_), .B(adder_bOperand_10_bF_buf3), .Y(divider_absoluteValue_B_flipSign_result_10_) );
	INVX1 INVX1_1512 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf2), .Y(_10911_) );
	AOI22X1 AOI22X1_245 ( .gnd(gnd), .vdd(vdd), .A(_10901_), .B(_10903_), .C(_10906_), .D(_10907_), .Y(_10912_) );
	NAND2X1 NAND2X1_1924 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf2), .B(_11054__bF_buf0), .Y(_10913_) );
	INVX1 INVX1_1513 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf1), .Y(_10914_) );
	NAND2X1 NAND2X1_1925 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf0), .B(_10914_), .Y(_10915_) );
	NAND2X1 NAND2X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .B(_10915_), .Y(_10916_) );
	NAND3X1 NAND3X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10916_), .C(_10900_), .Y(_10917_) );
	NAND2X1 NAND2X1_1927 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf1), .B(_11054__bF_buf4), .Y(_10918_) );
	NAND2X1 NAND2X1_1928 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(_10911_), .Y(_10919_) );
	NAND2X1 NAND2X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_10918_), .B(_10919_), .Y(_10920_) );
	NAND2X1 NAND2X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_10920_), .B(_10917_), .Y(_10921_) );
	OAI21X1 OAI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_10911_), .B(_10917_), .C(_10921_), .Y(divider_absoluteValue_B_flipSign_result_11_) );
	NAND2X1 NAND2X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10900_), .Y(_10922_) );
	AOI22X1 AOI22X1_246 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .B(_10915_), .C(_10918_), .D(_10919_), .Y(_10923_) );
	INVX1 INVX1_1514 ( .gnd(gnd), .vdd(vdd), .A(_10923_), .Y(_10924_) );
	OAI21X1 OAI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_10924_), .B(_10922_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf4), .Y(_10925_) );
	XNOR2X1 XNOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_10925_), .B(adder_bOperand_12_bF_buf2), .Y(divider_absoluteValue_B_flipSign_result_12_) );
	INVX1 INVX1_1515 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf3), .Y(_10926_) );
	NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_10924_), .B(_10922_), .Y(_10927_) );
	NAND2X1 NAND2X1_1932 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf1), .B(_11054__bF_buf3), .Y(_10928_) );
	INVX1 INVX1_1516 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf0), .Y(_10929_) );
	NAND2X1 NAND2X1_1933 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(_10929_), .Y(_10930_) );
	NAND2X1 NAND2X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_10928_), .B(_10930_), .Y(_10931_) );
	NAND2X1 NAND2X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_10931_), .B(_10927_), .Y(_10932_) );
	NAND2X1 NAND2X1_1936 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf2), .B(_11054__bF_buf2), .Y(_10933_) );
	NAND2X1 NAND2X1_1937 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf2), .B(_10926_), .Y(_10934_) );
	NAND2X1 NAND2X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_10933_), .B(_10934_), .Y(_10935_) );
	NAND2X1 NAND2X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_10935_), .B(_10932_), .Y(_10936_) );
	OAI21X1 OAI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_10926_), .B(_10932_), .C(_10936_), .Y(divider_absoluteValue_B_flipSign_result_13_) );
	INVX1 INVX1_1517 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf3), .Y(_10937_) );
	NAND3X1 NAND3X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10923_), .C(_10900_), .Y(_10938_) );
	AOI22X1 AOI22X1_247 ( .gnd(gnd), .vdd(vdd), .A(_10928_), .B(_10930_), .C(_10933_), .D(_10934_), .Y(_10939_) );
	INVX1 INVX1_1518 ( .gnd(gnd), .vdd(vdd), .A(_10939_), .Y(_10940_) );
	NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_10940_), .B(_10938_), .Y(_10941_) );
	NAND2X1 NAND2X1_1940 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf2), .B(_11054__bF_buf1), .Y(_10942_) );
	NAND2X1 NAND2X1_1941 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf1), .B(_10937_), .Y(_10943_) );
	NAND2X1 NAND2X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_10942_), .B(_10943_), .Y(_10944_) );
	AOI21X1 AOI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_10927_), .B(_10939_), .C(_10944_), .Y(_10945_) );
	AOI21X1 AOI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_10937_), .B(_10941_), .C(_10945_), .Y(divider_absoluteValue_B_flipSign_result_14_) );
	INVX1 INVX1_1519 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf3), .Y(_10946_) );
	NAND2X1 NAND2X1_1943 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf2), .B(_11054__bF_buf0), .Y(_10947_) );
	NAND2X1 NAND2X1_1944 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf0), .B(_10946_), .Y(_10948_) );
	NAND2X1 NAND2X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_10947_), .B(_10948_), .Y(_10949_) );
	INVX1 INVX1_1520 ( .gnd(gnd), .vdd(vdd), .A(_10949_), .Y(_10950_) );
	NAND2X1 NAND2X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_10944_), .B(_10941_), .Y(_10951_) );
	MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_10950_), .B(_10946_), .S(_10951_), .Y(divider_absoluteValue_B_flipSign_result_15_) );
	NAND2X1 NAND2X1_1947 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_bF_buf3), .B(_11054__bF_buf4), .Y(_10952_) );
	NAND2X1 NAND2X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10923_), .Y(_10953_) );
	AOI22X1 AOI22X1_248 ( .gnd(gnd), .vdd(vdd), .A(_10942_), .B(_10943_), .C(_10947_), .D(_10948_), .Y(_10954_) );
	NAND2X1 NAND2X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_10939_), .B(_10954_), .Y(_10955_) );
	NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(_10953_), .B(_10955_), .Y(_10956_) );
	AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_10956_), .B(_10900_), .Y(_10957_) );
	INVX1 INVX1_1521 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_bF_buf2), .Y(_10958_) );
	NAND2X1 NAND2X1_1950 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(_10958_), .Y(_10959_) );
	NAND2X1 NAND2X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_10952_), .B(_10959_), .Y(_10960_) );
	XNOR2X1 XNOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_10957_), .B(_10960_), .Y(_10961_) );
	OAI21X1 OAI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_11054__bF_buf3), .B(_10961_), .C(_10952_), .Y(divider_absoluteValue_B_flipSign_result_16_) );
	INVX1 INVX1_1522 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf3), .Y(_10962_) );
	NAND2X1 NAND2X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_10912_), .B(_10954_), .Y(_10963_) );
	NAND2X1 NAND2X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_10923_), .B(_10939_), .Y(_10964_) );
	NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(_10963_), .B(_10964_), .Y(_10965_) );
	AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_10965_), .B(_10900_), .Y(_10966_) );
	NAND2X1 NAND2X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_10960_), .B(_10966_), .Y(_10967_) );
	INVX1 INVX1_1523 ( .gnd(gnd), .vdd(vdd), .A(_10957_), .Y(_10968_) );
	INVX1 INVX1_1524 ( .gnd(gnd), .vdd(vdd), .A(_10960_), .Y(_10969_) );
	NAND2X1 NAND2X1_1955 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf2), .B(_11054__bF_buf2), .Y(_10970_) );
	NAND2X1 NAND2X1_1956 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf4), .B(_10962_), .Y(_10971_) );
	NAND2X1 NAND2X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_10970_), .B(_10971_), .Y(_10972_) );
	OAI21X1 OAI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_10969_), .B(_10968_), .C(_10972_), .Y(_10973_) );
	OAI21X1 OAI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_10962_), .B(_10967_), .C(_10973_), .Y(divider_absoluteValue_B_flipSign_result_17_) );
	INVX1 INVX1_1525 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf2), .Y(_10974_) );
	AOI22X1 AOI22X1_249 ( .gnd(gnd), .vdd(vdd), .A(_10952_), .B(_10959_), .C(_10970_), .D(_10971_), .Y(_10975_) );
	AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_10966_), .B(_10975_), .Y(_10976_) );
	NAND2X1 NAND2X1_1958 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf1), .B(_11054__bF_buf1), .Y(_10977_) );
	NAND2X1 NAND2X1_1959 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(_10974_), .Y(_10978_) );
	NAND2X1 NAND2X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_10977_), .B(_10978_), .Y(_10979_) );
	NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_10979_), .B(_10976_), .Y(_10980_) );
	AOI21X1 AOI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_10974_), .B(_10976_), .C(_10980_), .Y(divider_absoluteValue_B_flipSign_result_18_) );
	INVX1 INVX1_1526 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf1), .Y(_10981_) );
	NAND2X1 NAND2X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_10979_), .B(_10976_), .Y(_10982_) );
	XOR2X1 XOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf2), .B(adder_bOperand_19_bF_buf0), .Y(_10983_) );
	NAND2X1 NAND2X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_10983_), .B(_10982_), .Y(_10984_) );
	OAI21X1 OAI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_10981_), .B(_10982_), .C(_10984_), .Y(divider_absoluteValue_B_flipSign_result_19_) );
	NAND3X1 NAND3X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_10979_), .B(_10983_), .C(_10975_), .Y(_10985_) );
	OAI21X1 OAI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_10985_), .B(_10968_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf1), .Y(_10986_) );
	XNOR2X1 XNOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_10986_), .B(adder_bOperand_20_bF_buf0), .Y(divider_absoluteValue_B_flipSign_result_20_) );
	INVX1 INVX1_1527 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf2), .Y(_10987_) );
	NAND2X1 NAND2X1_1963 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf1), .B(_11054__bF_buf0), .Y(_10988_) );
	NAND2X1 NAND2X1_1964 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf0), .B(_10987_), .Y(_10989_) );
	AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_10988_), .B(_10989_), .Y(_10990_) );
	INVX1 INVX1_1528 ( .gnd(gnd), .vdd(vdd), .A(_10985_), .Y(_10991_) );
	NAND2X1 NAND2X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_10991_), .B(_10966_), .Y(_10992_) );
	NAND2X1 NAND2X1_1966 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf3), .B(_11054__bF_buf4), .Y(_10993_) );
	INVX1 INVX1_1529 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf2), .Y(_10994_) );
	NAND2X1 NAND2X1_1967 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(_10994_), .Y(_10995_) );
	AOI21X1 AOI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_10993_), .B(_10995_), .C(_10992_), .Y(_10996_) );
	MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_10987_), .B(_10990_), .S(_10996_), .Y(divider_absoluteValue_B_flipSign_result_21_) );
	INVX1 INVX1_1530 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf2), .Y(_10997_) );
	NAND2X1 NAND2X1_1968 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf1), .B(_11054__bF_buf3), .Y(_10998_) );
	NAND2X1 NAND2X1_1969 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf4), .B(_10997_), .Y(_10999_) );
	NAND2X1 NAND2X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_10998_), .B(_10999_), .Y(_11000_) );
	INVX1 INVX1_1531 ( .gnd(gnd), .vdd(vdd), .A(_11000_), .Y(_11001_) );
	AOI22X1 AOI22X1_250 ( .gnd(gnd), .vdd(vdd), .A(_10993_), .B(_10995_), .C(_10988_), .D(_10989_), .Y(_11002_) );
	INVX1 INVX1_1532 ( .gnd(gnd), .vdd(vdd), .A(_11002_), .Y(_11003_) );
	NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_11003_), .B(_10992_), .Y(_11004_) );
	MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_10997_), .B(_11001_), .S(_11004_), .Y(divider_absoluteValue_B_flipSign_result_22_) );
	XOR2X1 XOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(adder_bOperand_23_), .Y(_11005_) );
	INVX1 INVX1_1533 ( .gnd(gnd), .vdd(vdd), .A(_11005_), .Y(_11006_) );
	NAND2X1 NAND2X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_10991_), .B(_10957_), .Y(_11007_) );
	NOR3X1 NOR3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_11001_), .B(_11003_), .C(_11007_), .Y(_11008_) );
	NAND3X1 NAND3X1_2276 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_23_), .B(_11000_), .C(_11004_), .Y(_11009_) );
	OAI21X1 OAI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_11006_), .B(_11008_), .C(_11009_), .Y(divider_absoluteValue_B_flipSign_result_23_) );
	NAND2X1 NAND2X1_1972 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .B(_11054__bF_buf2), .Y(_11010_) );
	INVX1 INVX1_1534 ( .gnd(gnd), .vdd(vdd), .A(_11010_), .Y(_11011_) );
	NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .B(_11054__bF_buf1), .Y(_11012_) );
	OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_11011_), .B(_11012_), .Y(_11013_) );
	NAND3X1 NAND3X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_11000_), .B(_11005_), .C(_11002_), .Y(_11014_) );
	NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_10985_), .B(_11014_), .Y(_11015_) );
	NAND3X1 NAND3X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_10900_), .B(_10956_), .C(_11015_), .Y(_11016_) );
	XOR2X1 XOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_11016_), .B(_11013_), .Y(_11017_) );
	OAI21X1 OAI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_11054__bF_buf0), .B(_11017_), .C(_11010_), .Y(divider_absoluteValue_B_flipSign_result_24_) );
	OAI21X1 OAI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .B(_11016_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf2), .Y(_11018_) );
	XNOR2X1 XNOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_11018_), .B(adder_bOperand_25_), .Y(divider_absoluteValue_B_flipSign_result_25_) );
	XOR2X1 XOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf1), .B(adder_bOperand_25_), .Y(_11019_) );
	OAI21X1 OAI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_11012_), .B(_11011_), .C(_11019_), .Y(_11020_) );
	OAI21X1 OAI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .B(_11016_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf0), .Y(_11021_) );
	XNOR2X1 XNOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_11021_), .B(adder_bOperand_26_), .Y(divider_absoluteValue_B_flipSign_result_26_) );
	XOR2X1 XOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(adder_bOperand_27_), .Y(_11022_) );
	INVX1 INVX1_1535 ( .gnd(gnd), .vdd(vdd), .A(_11022_), .Y(_11023_) );
	NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .B(_11016_), .Y(_11024_) );
	XOR2X1 XOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf4), .B(adder_bOperand_26_), .Y(_11025_) );
	NAND2X1 NAND2X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_11025_), .B(_11024_), .Y(_11026_) );
	NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_27_), .B(_11026_), .Y(_11027_) );
	AOI21X1 AOI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_11023_), .B(_11026_), .C(_11027_), .Y(divider_absoluteValue_B_flipSign_result_27_) );
	INVX1 INVX1_1536 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .Y(_11028_) );
	AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_11025_), .B(_11022_), .Y(_11029_) );
	NAND2X1 NAND2X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_11029_), .B(_11028_), .Y(_11030_) );
	OAI21X1 OAI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_11030_), .B(_11016_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf3), .Y(_11031_) );
	XNOR2X1 XNOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_11031_), .B(adder_bOperand_28_), .Y(divider_absoluteValue_B_flipSign_result_28_) );
	XOR2X1 XOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf2), .B(adder_bOperand_29_), .Y(_11032_) );
	INVX1 INVX1_1537 ( .gnd(gnd), .vdd(vdd), .A(_11032_), .Y(_11033_) );
	NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_11030_), .B(_11016_), .Y(_11034_) );
	XNOR2X1 XNOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf1), .B(adder_bOperand_28_), .Y(_11035_) );
	INVX1 INVX1_1538 ( .gnd(gnd), .vdd(vdd), .A(_11035_), .Y(_11036_) );
	NAND2X1 NAND2X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_11036_), .B(_11034_), .Y(_11037_) );
	NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_29_), .B(_11037_), .Y(_11038_) );
	AOI21X1 AOI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_11033_), .B(_11037_), .C(_11038_), .Y(divider_absoluteValue_B_flipSign_result_29_) );
	INVX1 INVX1_1539 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_30_), .Y(_11039_) );
	NAND2X1 NAND2X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_11032_), .B(_11036_), .Y(_11040_) );
	NOR3X1 NOR3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_11030_), .B(_11040_), .C(_11016_), .Y(_11041_) );
	OAI21X1 OAI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_11054__bF_buf4), .B(_11041_), .C(_11039_), .Y(_11042_) );
	INVX1 INVX1_1540 ( .gnd(gnd), .vdd(vdd), .A(_11040_), .Y(_11043_) );
	NAND2X1 NAND2X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_11043_), .B(_11034_), .Y(_11044_) );
	NAND3X1 NAND3X1_2279 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf0), .B(adder_bOperand_30_), .C(_11044_), .Y(_11045_) );
	AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_11045_), .B(_11042_), .Y(divider_absoluteValue_B_flipSign_result_30_) );
	INVX1 INVX1_1541 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_msb), .Y(_11046_) );
	NAND3X1 NAND3X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_11039_), .B(_11043_), .C(_11034_), .Y(_11047_) );
	NAND3X1 NAND3X1_2281 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf5), .B(_11046_), .C(_11047_), .Y(_11048_) );
	INVX1 INVX1_1542 ( .gnd(gnd), .vdd(vdd), .A(_11030_), .Y(_11049_) );
	NAND3X1 NAND3X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_11015_), .B(_11049_), .C(_10957_), .Y(_11050_) );
	OAI21X1 OAI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_11040_), .B(_11050_), .C(divider_absoluteValue_B_flipSign_flip_bF_buf4), .Y(_11051_) );
	NAND2X1 NAND2X1_1978 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_flipSign_flip_bF_buf3), .B(adder_bOperand_30_), .Y(_11052_) );
	NAND3X1 NAND3X1_2283 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_msb), .B(_11052_), .C(_11051_), .Y(_11053_) );
	NAND2X1 NAND2X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_11048_), .B(_11053_), .Y(divider_absoluteValue_B_flipSign_result_31_) );
	BUFX4 BUFX4_1976 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .Y(divider_absoluteValue_B_flipSign_result_0_) );
	INVX8 INVX8_43 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf5), .Y(_11252_) );
	NAND2X1 NAND2X1_1980 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_1_bF_buf3), .B(_11252__bF_buf4), .Y(_11253_) );
	XOR2X1 XOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(divider_divuResult_0_bF_buf4), .Y(_11254_) );
	XOR2X1 XOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf3), .B(divider_divuResult_1_bF_buf2), .Y(_11255_) );
	NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_11254_), .B(_11255_), .Y(_11256_) );
	OAI21X1 OAI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf3), .B(divider_divuResult_1_bF_buf1), .C(divider_divFlip_bF_buf2), .Y(_11257_) );
	OAI21X1 OAI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_11257_), .B(_11256_), .C(_11253_), .Y(divideOut_1_) );
	INVX1 INVX1_1543 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf2), .Y(_11258_) );
	AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_11254_), .B(_11255_), .Y(_11259_) );
	INVX1 INVX1_1544 ( .gnd(gnd), .vdd(vdd), .A(_11259_), .Y(_11260_) );
	OAI21X1 OAI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf1), .B(_11260_), .C(divider_divFlip_bF_buf1), .Y(_11261_) );
	NOR2X1 NOR2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_11258_), .B(_11259_), .Y(_11262_) );
	OAI22X1 OAI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(_11258_), .C(_11262_), .D(_11261_), .Y(divideOut_2_) );
	XNOR2X1 XNOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_11261_), .B(divider_divuResult_3_bF_buf0), .Y(divideOut_3_) );
	NAND2X1 NAND2X1_1981 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf0), .B(_11252__bF_buf3), .Y(_11263_) );
	NAND3X1 NAND3X1_2284 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_2_bF_buf0), .B(divider_divuResult_3_bF_buf7), .C(_11252__bF_buf2), .Y(_11264_) );
	INVX1 INVX1_1545 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_3_bF_buf6), .Y(_11265_) );
	NAND3X1 NAND3X1_2285 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf5), .B(_11258_), .C(_11265_), .Y(_11266_) );
	NAND2X1 NAND2X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_11264_), .B(_11266_), .Y(_11267_) );
	NAND3X1 NAND3X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_11254_), .B(_11255_), .C(_11267_), .Y(_11268_) );
	INVX1 INVX1_1546 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_4_bF_buf6), .Y(_11269_) );
	NAND2X1 NAND2X1_1983 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(_11269_), .Y(_11270_) );
	NAND2X1 NAND2X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_11263_), .B(_11270_), .Y(_11271_) );
	XOR2X1 XOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_11268_), .B(_11271_), .Y(_11272_) );
	OAI21X1 OAI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_11252__bF_buf1), .B(_11272_), .C(_11263_), .Y(divideOut_4_) );
	INVX1 INVX1_1547 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf2), .Y(_11273_) );
	NAND3X1 NAND3X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_11267_), .B(_11271_), .C(_11259_), .Y(_11274_) );
	NAND2X1 NAND2X1_1985 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf1), .B(_11252__bF_buf0), .Y(_11275_) );
	NAND2X1 NAND2X1_1986 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf3), .B(_11273_), .Y(_11276_) );
	NAND2X1 NAND2X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11276_), .Y(_11277_) );
	NAND2X1 NAND2X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_11277_), .B(_11274_), .Y(_11278_) );
	OAI21X1 OAI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_11273_), .B(_11274_), .C(_11278_), .Y(divideOut_5_) );
	OAI21X1 OAI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_5_bF_buf0), .B(_11274_), .C(divider_divFlip_bF_buf2), .Y(_11279_) );
	XNOR2X1 XNOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_11279_), .B(divider_divuResult_6_bF_buf0), .Y(divideOut_6_) );
	INVX1 INVX1_1548 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf1), .Y(_11082_) );
	AOI21X1 AOI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_11275_), .B(_11276_), .C(_11274_), .Y(_11083_) );
	NAND2X1 NAND2X1_1989 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf6), .B(_11252__bF_buf4), .Y(_11084_) );
	INVX1 INVX1_1549 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_6_bF_buf5), .Y(_11085_) );
	NAND2X1 NAND2X1_1990 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf1), .B(_11085_), .Y(_11086_) );
	NAND2X1 NAND2X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_11084_), .B(_11086_), .Y(_11087_) );
	NAND2X1 NAND2X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .B(_11083_), .Y(_11088_) );
	NAND2X1 NAND2X1_1993 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_7_bF_buf0), .B(_11252__bF_buf3), .Y(_11089_) );
	NAND2X1 NAND2X1_1994 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(_11082_), .Y(_11090_) );
	NAND2X1 NAND2X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_11089_), .B(_11090_), .Y(_11091_) );
	NAND2X1 NAND2X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_11091_), .B(_11088_), .Y(_11092_) );
	OAI21X1 OAI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_11082_), .B(_11088_), .C(_11092_), .Y(divideOut_7_) );
	AOI22X1 AOI22X1_251 ( .gnd(gnd), .vdd(vdd), .A(_11263_), .B(_11270_), .C(_11275_), .D(_11276_), .Y(_11093_) );
	AOI22X1 AOI22X1_252 ( .gnd(gnd), .vdd(vdd), .A(_11084_), .B(_11086_), .C(_11089_), .D(_11090_), .Y(_11094_) );
	NAND2X1 NAND2X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_11093_), .B(_11094_), .Y(_11095_) );
	OAI21X1 OAI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_11268_), .B(_11095_), .C(divider_divFlip_bF_buf5), .Y(_11096_) );
	XNOR2X1 XNOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_11096_), .B(divider_divuResult_8_bF_buf1), .Y(divideOut_8_) );
	INVX1 INVX1_1550 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf1), .Y(_11097_) );
	NOR2X1 NOR2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_11268_), .B(_11095_), .Y(_11098_) );
	NAND2X1 NAND2X1_1998 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf0), .B(_11252__bF_buf2), .Y(_11099_) );
	INVX1 INVX1_1551 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_8_bF_buf6), .Y(_11100_) );
	NAND2X1 NAND2X1_1999 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(_11100_), .Y(_11101_) );
	NAND2X1 NAND2X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_11099_), .B(_11101_), .Y(_11102_) );
	NAND2X1 NAND2X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_11102_), .B(_11098_), .Y(_11103_) );
	NAND2X1 NAND2X1_2002 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf0), .B(_11252__bF_buf1), .Y(_11104_) );
	NAND2X1 NAND2X1_2003 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf3), .B(_11097_), .Y(_11105_) );
	NAND2X1 NAND2X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_11104_), .B(_11105_), .Y(_11106_) );
	NAND2X1 NAND2X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_11106_), .B(_11103_), .Y(_11107_) );
	OAI21X1 OAI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_11097_), .B(_11103_), .C(_11107_), .Y(divideOut_9_) );
	OAI21X1 OAI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_9_bF_buf5), .B(_11103_), .C(divider_divFlip_bF_buf2), .Y(_11108_) );
	XNOR2X1 XNOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_11108_), .B(divider_divuResult_10_bF_buf2), .Y(divideOut_10_) );
	INVX1 INVX1_1552 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf2), .Y(_11109_) );
	AOI22X1 AOI22X1_253 ( .gnd(gnd), .vdd(vdd), .A(_11099_), .B(_11101_), .C(_11104_), .D(_11105_), .Y(_11110_) );
	NAND2X1 NAND2X1_2006 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf1), .B(_11252__bF_buf0), .Y(_11111_) );
	INVX1 INVX1_1553 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_10_bF_buf0), .Y(_11112_) );
	NAND2X1 NAND2X1_2007 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf1), .B(_11112_), .Y(_11113_) );
	NAND2X1 NAND2X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_11111_), .B(_11113_), .Y(_11114_) );
	NAND3X1 NAND3X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11114_), .C(_11098_), .Y(_11115_) );
	NAND2X1 NAND2X1_2009 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_11_bF_buf1), .B(_11252__bF_buf4), .Y(_11116_) );
	NAND2X1 NAND2X1_2010 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(_11109_), .Y(_11117_) );
	NAND2X1 NAND2X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_11116_), .B(_11117_), .Y(_11118_) );
	NAND2X1 NAND2X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_11118_), .B(_11115_), .Y(_11119_) );
	OAI21X1 OAI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_11109_), .B(_11115_), .C(_11119_), .Y(divideOut_11_) );
	NAND2X1 NAND2X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11098_), .Y(_11120_) );
	AOI22X1 AOI22X1_254 ( .gnd(gnd), .vdd(vdd), .A(_11111_), .B(_11113_), .C(_11116_), .D(_11117_), .Y(_11121_) );
	INVX1 INVX1_1554 ( .gnd(gnd), .vdd(vdd), .A(_11121_), .Y(_11122_) );
	OAI21X1 OAI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_11122_), .B(_11120_), .C(divider_divFlip_bF_buf5), .Y(_11123_) );
	XNOR2X1 XNOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_11123_), .B(divider_divuResult_12_bF_buf4), .Y(divideOut_12_) );
	INVX1 INVX1_1555 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf5), .Y(_11124_) );
	NOR2X1 NOR2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_11122_), .B(_11120_), .Y(_11125_) );
	NAND2X1 NAND2X1_2014 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf3), .B(_11252__bF_buf3), .Y(_11126_) );
	INVX1 INVX1_1556 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_12_bF_buf2), .Y(_11127_) );
	NAND2X1 NAND2X1_2015 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(_11127_), .Y(_11128_) );
	NAND2X1 NAND2X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_11126_), .B(_11128_), .Y(_11129_) );
	NAND2X1 NAND2X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_11129_), .B(_11125_), .Y(_11130_) );
	NAND2X1 NAND2X1_2018 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_13_bF_buf4), .B(_11252__bF_buf2), .Y(_11131_) );
	NAND2X1 NAND2X1_2019 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf3), .B(_11124_), .Y(_11132_) );
	NAND2X1 NAND2X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_11131_), .B(_11132_), .Y(_11133_) );
	NAND2X1 NAND2X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_11133_), .B(_11130_), .Y(_11134_) );
	OAI21X1 OAI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_11124_), .B(_11130_), .C(_11134_), .Y(divideOut_13_) );
	INVX1 INVX1_1557 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf1), .Y(_11135_) );
	NAND3X1 NAND3X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11121_), .C(_11098_), .Y(_11136_) );
	AOI22X1 AOI22X1_255 ( .gnd(gnd), .vdd(vdd), .A(_11126_), .B(_11128_), .C(_11131_), .D(_11132_), .Y(_11137_) );
	INVX1 INVX1_1558 ( .gnd(gnd), .vdd(vdd), .A(_11137_), .Y(_11138_) );
	NOR2X1 NOR2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11136_), .Y(_11139_) );
	NAND2X1 NAND2X1_2022 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_14_bF_buf0), .B(_11252__bF_buf1), .Y(_11140_) );
	NAND2X1 NAND2X1_2023 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf2), .B(_11135_), .Y(_11141_) );
	NAND2X1 NAND2X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_11140_), .B(_11141_), .Y(_11142_) );
	AOI21X1 AOI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_11125_), .B(_11137_), .C(_11142_), .Y(_11143_) );
	AOI21X1 AOI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_11135_), .B(_11139_), .C(_11143_), .Y(divideOut_14_) );
	INVX1 INVX1_1559 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf4), .Y(_11144_) );
	NAND2X1 NAND2X1_2025 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_15_bF_buf3), .B(_11252__bF_buf0), .Y(_11145_) );
	NAND2X1 NAND2X1_2026 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf1), .B(_11144_), .Y(_11146_) );
	NAND2X1 NAND2X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_11145_), .B(_11146_), .Y(_11147_) );
	INVX1 INVX1_1560 ( .gnd(gnd), .vdd(vdd), .A(_11147_), .Y(_11148_) );
	NAND2X1 NAND2X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_11142_), .B(_11139_), .Y(_11149_) );
	MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_11148_), .B(_11144_), .S(_11149_), .Y(divideOut_15_) );
	NAND2X1 NAND2X1_2029 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf5), .B(_11252__bF_buf4), .Y(_11150_) );
	NAND2X1 NAND2X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11121_), .Y(_11151_) );
	AOI22X1 AOI22X1_256 ( .gnd(gnd), .vdd(vdd), .A(_11140_), .B(_11141_), .C(_11145_), .D(_11146_), .Y(_11152_) );
	NAND2X1 NAND2X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_11137_), .B(_11152_), .Y(_11153_) );
	NOR2X1 NOR2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_11151_), .B(_11153_), .Y(_11154_) );
	AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_11154_), .B(_11098_), .Y(_11155_) );
	INVX1 INVX1_1561 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_16_bF_buf4), .Y(_11156_) );
	NAND2X1 NAND2X1_2032 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(_11156_), .Y(_11157_) );
	NAND2X1 NAND2X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_11150_), .B(_11157_), .Y(_11158_) );
	XNOR2X1 XNOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(_11158_), .Y(_11159_) );
	OAI21X1 OAI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_11252__bF_buf3), .B(_11159_), .C(_11150_), .Y(divideOut_16_) );
	INVX1 INVX1_1562 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_17_bF_buf1), .Y(_11160_) );
	NAND2X1 NAND2X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_11110_), .B(_11152_), .Y(_11161_) );
	NAND2X1 NAND2X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_11121_), .B(_11137_), .Y(_11162_) );
	NOR2X1 NOR2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_11161_), .B(_11162_), .Y(_11163_) );
	AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_11163_), .B(_11098_), .Y(_11164_) );
	NAND2X1 NAND2X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .B(_11164_), .Y(_11165_) );
	INVX1 INVX1_1563 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .Y(_11166_) );
	INVX1 INVX1_1564 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .Y(_11167_) );
	NAND2X1 NAND2X1_2037 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_17_bF_buf0), .B(_11252__bF_buf2), .Y(_11168_) );
	NAND2X1 NAND2X1_2038 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf5), .B(_11160_), .Y(_11169_) );
	NAND2X1 NAND2X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_11168_), .B(_11169_), .Y(_11170_) );
	OAI21X1 OAI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_11167_), .B(_11166_), .C(_11170_), .Y(_11171_) );
	OAI21X1 OAI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_11160_), .B(_11165_), .C(_11171_), .Y(divideOut_17_) );
	INVX1 INVX1_1565 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf0), .Y(_11172_) );
	AOI22X1 AOI22X1_257 ( .gnd(gnd), .vdd(vdd), .A(_11150_), .B(_11157_), .C(_11168_), .D(_11169_), .Y(_11173_) );
	AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_11164_), .B(_11173_), .Y(_11174_) );
	NAND2X1 NAND2X1_2040 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_18_bF_buf5), .B(_11252__bF_buf1), .Y(_11175_) );
	NAND2X1 NAND2X1_2041 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(_11172_), .Y(_11176_) );
	NAND2X1 NAND2X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_11175_), .B(_11176_), .Y(_11177_) );
	NOR2X1 NOR2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_11177_), .B(_11174_), .Y(_11178_) );
	AOI21X1 AOI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_11172_), .B(_11174_), .C(_11178_), .Y(divideOut_18_) );
	INVX1 INVX1_1566 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_19_bF_buf4), .Y(_11179_) );
	NAND2X1 NAND2X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_11177_), .B(_11174_), .Y(_11180_) );
	XOR2X1 XOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf3), .B(divider_divuResult_19_bF_buf3), .Y(_11181_) );
	NAND2X1 NAND2X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_11181_), .B(_11180_), .Y(_11182_) );
	OAI21X1 OAI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_11179_), .B(_11180_), .C(_11182_), .Y(divideOut_19_) );
	NAND3X1 NAND3X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_11177_), .B(_11181_), .C(_11173_), .Y(_11183_) );
	OAI21X1 OAI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_11183_), .B(_11166_), .C(divider_divFlip_bF_buf2), .Y(_11184_) );
	XNOR2X1 XNOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_11184_), .B(divider_divuResult_20_bF_buf3), .Y(divideOut_20_) );
	INVX1 INVX1_1567 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_bF_buf3), .Y(_11185_) );
	NAND2X1 NAND2X1_2045 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_21_bF_buf2), .B(_11252__bF_buf0), .Y(_11186_) );
	NAND2X1 NAND2X1_2046 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf1), .B(_11185_), .Y(_11187_) );
	AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_11186_), .B(_11187_), .Y(_11188_) );
	INVX1 INVX1_1568 ( .gnd(gnd), .vdd(vdd), .A(_11183_), .Y(_11189_) );
	NAND2X1 NAND2X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_11189_), .B(_11164_), .Y(_11190_) );
	NAND2X1 NAND2X1_2048 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf2), .B(_11252__bF_buf4), .Y(_11191_) );
	INVX1 INVX1_1569 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_20_bF_buf1), .Y(_11192_) );
	NAND2X1 NAND2X1_2049 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(_11192_), .Y(_11193_) );
	AOI21X1 AOI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_11191_), .B(_11193_), .C(_11190_), .Y(_11194_) );
	MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_11185_), .B(_11188_), .S(_11194_), .Y(divideOut_21_) );
	INVX1 INVX1_1570 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_22_), .Y(_11195_) );
	NAND2X1 NAND2X1_2050 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_22_), .B(_11252__bF_buf3), .Y(_11196_) );
	NAND2X1 NAND2X1_2051 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf5), .B(_11195_), .Y(_11197_) );
	NAND2X1 NAND2X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_11196_), .B(_11197_), .Y(_11198_) );
	INVX1 INVX1_1571 ( .gnd(gnd), .vdd(vdd), .A(_11198_), .Y(_11199_) );
	AOI22X1 AOI22X1_258 ( .gnd(gnd), .vdd(vdd), .A(_11191_), .B(_11193_), .C(_11186_), .D(_11187_), .Y(_11200_) );
	INVX1 INVX1_1572 ( .gnd(gnd), .vdd(vdd), .A(_11200_), .Y(_11201_) );
	NOR2X1 NOR2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_11201_), .B(_11190_), .Y(_11202_) );
	MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_11195_), .B(_11199_), .S(_11202_), .Y(divideOut_22_) );
	XOR2X1 XOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(divider_divuResult_23_), .Y(_11203_) );
	INVX1 INVX1_1573 ( .gnd(gnd), .vdd(vdd), .A(_11203_), .Y(_11204_) );
	NAND2X1 NAND2X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_11189_), .B(_11155_), .Y(_11205_) );
	NOR3X1 NOR3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_11199_), .B(_11201_), .C(_11205_), .Y(_11206_) );
	NAND3X1 NAND3X1_2291 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_23_), .B(_11198_), .C(_11202_), .Y(_11207_) );
	OAI21X1 OAI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_11204_), .B(_11206_), .C(_11207_), .Y(divideOut_23_) );
	NAND2X1 NAND2X1_2054 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf2), .B(_11252__bF_buf2), .Y(_11208_) );
	INVX1 INVX1_1574 ( .gnd(gnd), .vdd(vdd), .A(_11208_), .Y(_11209_) );
	NOR2X1 NOR2X1_730 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf1), .B(_11252__bF_buf1), .Y(_11210_) );
	OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_11209_), .B(_11210_), .Y(_11211_) );
	NAND3X1 NAND3X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_11198_), .B(_11203_), .C(_11200_), .Y(_11212_) );
	NOR2X1 NOR2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_11183_), .B(_11212_), .Y(_11213_) );
	NAND3X1 NAND3X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_11098_), .B(_11154_), .C(_11213_), .Y(_11214_) );
	XOR2X1 XOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_11214_), .B(_11211_), .Y(_11215_) );
	OAI21X1 OAI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_11252__bF_buf0), .B(_11215_), .C(_11208_), .Y(divideOut_24_) );
	OAI21X1 OAI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_24_bF_buf0), .B(_11214_), .C(divider_divFlip_bF_buf3), .Y(_11216_) );
	XNOR2X1 XNOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_11216_), .B(divider_divuResult_25_), .Y(divideOut_25_) );
	XOR2X1 XOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf2), .B(divider_divuResult_25_), .Y(_11217_) );
	OAI21X1 OAI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_11210_), .B(_11209_), .C(_11217_), .Y(_11218_) );
	OAI21X1 OAI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_11218_), .B(_11214_), .C(divider_divFlip_bF_buf1), .Y(_11219_) );
	XNOR2X1 XNOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_11219_), .B(divider_divuResult_26_), .Y(divideOut_26_) );
	XOR2X1 XOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(divider_divuResult_27_), .Y(_11220_) );
	INVX1 INVX1_1575 ( .gnd(gnd), .vdd(vdd), .A(_11220_), .Y(_11221_) );
	NOR2X1 NOR2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_11218_), .B(_11214_), .Y(_11222_) );
	XOR2X1 XOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf5), .B(divider_divuResult_26_), .Y(_11223_) );
	NAND2X1 NAND2X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_11223_), .B(_11222_), .Y(_11224_) );
	NOR2X1 NOR2X1_733 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_27_), .B(_11224_), .Y(_11225_) );
	AOI21X1 AOI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_11221_), .B(_11224_), .C(_11225_), .Y(divideOut_27_) );
	INVX1 INVX1_1576 ( .gnd(gnd), .vdd(vdd), .A(_11218_), .Y(_11226_) );
	AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_11223_), .B(_11220_), .Y(_11227_) );
	NAND2X1 NAND2X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_11227_), .B(_11226_), .Y(_11228_) );
	OAI21X1 OAI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_11228_), .B(_11214_), .C(divider_divFlip_bF_buf4), .Y(_11229_) );
	XNOR2X1 XNOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_11229_), .B(divider_divuResult_28_), .Y(divideOut_28_) );
	XOR2X1 XOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf3), .B(divider_divuResult_29_), .Y(_11230_) );
	INVX1 INVX1_1577 ( .gnd(gnd), .vdd(vdd), .A(_11230_), .Y(_11231_) );
	NOR2X1 NOR2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_11228_), .B(_11214_), .Y(_11232_) );
	XNOR2X1 XNOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf2), .B(divider_divuResult_28_), .Y(_11233_) );
	INVX1 INVX1_1578 ( .gnd(gnd), .vdd(vdd), .A(_11233_), .Y(_11234_) );
	NAND2X1 NAND2X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_11234_), .B(_11232_), .Y(_11235_) );
	NOR2X1 NOR2X1_735 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_29_), .B(_11235_), .Y(_11236_) );
	AOI21X1 AOI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_11231_), .B(_11235_), .C(_11236_), .Y(divideOut_29_) );
	INVX1 INVX1_1579 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_30_), .Y(_11237_) );
	NAND2X1 NAND2X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_11230_), .B(_11234_), .Y(_11238_) );
	NOR3X1 NOR3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_11228_), .B(_11238_), .C(_11214_), .Y(_11239_) );
	OAI21X1 OAI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_11252__bF_buf4), .B(_11239_), .C(_11237_), .Y(_11240_) );
	INVX1 INVX1_1580 ( .gnd(gnd), .vdd(vdd), .A(_11238_), .Y(_11241_) );
	NAND2X1 NAND2X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_11241_), .B(_11232_), .Y(_11242_) );
	NAND3X1 NAND3X1_2294 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf1), .B(divider_divuResult_30_), .C(_11242_), .Y(_11243_) );
	AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_11243_), .B(_11240_), .Y(divideOut_30_) );
	INVX1 INVX1_1581 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_31_), .Y(_11244_) );
	NAND3X1 NAND3X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_11237_), .B(_11241_), .C(_11232_), .Y(_11245_) );
	NAND3X1 NAND3X1_2296 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf0), .B(_11244_), .C(_11245_), .Y(_11246_) );
	INVX1 INVX1_1582 ( .gnd(gnd), .vdd(vdd), .A(_11228_), .Y(_11247_) );
	NAND3X1 NAND3X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_11213_), .B(_11247_), .C(_11155_), .Y(_11248_) );
	OAI21X1 OAI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_11238_), .B(_11248_), .C(divider_divFlip_bF_buf5), .Y(_11249_) );
	NAND2X1 NAND2X1_2060 ( .gnd(gnd), .vdd(vdd), .A(divider_divFlip_bF_buf4), .B(divider_divuResult_30_), .Y(_11250_) );
	NAND3X1 NAND3X1_2298 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_31_), .B(_11250_), .C(_11249_), .Y(_11251_) );
	NAND2X1 NAND2X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_11246_), .B(_11251_), .Y(divideOut_31_) );
	BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(divider_divuResult_0_bF_buf2), .Y(divideOut_0_) );
	INVX8 INVX8_44 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf8), .Y(_11450_) );
	NAND2X1 NAND2X1_2062 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_1_), .B(_11450__bF_buf4), .Y(_11451_) );
	XOR2X1 XOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf7), .B(divider_flipSign_rem_operand_0_), .Y(_11452_) );
	XOR2X1 XOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(divider_flipSign_rem_operand_1_), .Y(_11453_) );
	NOR2X1 NOR2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_11452_), .B(_11453_), .Y(_11454_) );
	OAI21X1 OAI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_0_), .B(divider_flipSign_rem_operand_1_), .C(divider_a_isNegative_bF_buf5), .Y(_11455_) );
	OAI21X1 OAI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_11455_), .B(_11454_), .C(_11451_), .Y(divider_flipSign_rem_result_1_) );
	INVX1 INVX1_1583 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_2_), .Y(_11456_) );
	AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_11452_), .B(_11453_), .Y(_11457_) );
	INVX1 INVX1_1584 ( .gnd(gnd), .vdd(vdd), .A(_11457_), .Y(_11458_) );
	OAI21X1 OAI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_2_), .B(_11458_), .C(divider_a_isNegative_bF_buf4), .Y(_11459_) );
	NOR2X1 NOR2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_11456_), .B(_11457_), .Y(_11460_) );
	OAI22X1 OAI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(_11456_), .C(_11460_), .D(_11459_), .Y(divider_flipSign_rem_result_2_) );
	XNOR2X1 XNOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_11459_), .B(divider_flipSign_rem_operand_3_), .Y(divider_flipSign_rem_result_3_) );
	NAND2X1 NAND2X1_2063 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_4_), .B(_11450__bF_buf3), .Y(_11461_) );
	NAND3X1 NAND3X1_2299 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_2_), .B(divider_flipSign_rem_operand_3_), .C(_11450__bF_buf2), .Y(_11462_) );
	INVX1 INVX1_1585 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_3_), .Y(_11463_) );
	NAND3X1 NAND3X1_2300 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(_11456_), .C(_11463_), .Y(_11464_) );
	NAND2X1 NAND2X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_11462_), .B(_11464_), .Y(_11465_) );
	NAND3X1 NAND3X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_11452_), .B(_11453_), .C(_11465_), .Y(_11466_) );
	INVX1 INVX1_1586 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_4_), .Y(_11467_) );
	NAND2X1 NAND2X1_2065 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(_11467_), .Y(_11468_) );
	NAND2X1 NAND2X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_11461_), .B(_11468_), .Y(_11469_) );
	XOR2X1 XOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_11466_), .B(_11469_), .Y(_11470_) );
	OAI21X1 OAI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_11450__bF_buf1), .B(_11470_), .C(_11461_), .Y(divider_flipSign_rem_result_4_) );
	INVX1 INVX1_1587 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_5_), .Y(_11471_) );
	NAND3X1 NAND3X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_11465_), .B(_11469_), .C(_11457_), .Y(_11472_) );
	NAND2X1 NAND2X1_2067 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_5_), .B(_11450__bF_buf0), .Y(_11473_) );
	NAND2X1 NAND2X1_2068 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(_11471_), .Y(_11474_) );
	NAND2X1 NAND2X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_11473_), .B(_11474_), .Y(_11475_) );
	NAND2X1 NAND2X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_11475_), .B(_11472_), .Y(_11476_) );
	OAI21X1 OAI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_11471_), .B(_11472_), .C(_11476_), .Y(divider_flipSign_rem_result_5_) );
	OAI21X1 OAI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_5_), .B(_11472_), .C(divider_a_isNegative_bF_buf8), .Y(_11477_) );
	XNOR2X1 XNOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_11477_), .B(divider_flipSign_rem_operand_6_), .Y(divider_flipSign_rem_result_6_) );
	INVX1 INVX1_1588 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_7_), .Y(_11280_) );
	AOI21X1 AOI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_11473_), .B(_11474_), .C(_11472_), .Y(_11281_) );
	NAND2X1 NAND2X1_2071 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_6_), .B(_11450__bF_buf4), .Y(_11282_) );
	INVX1 INVX1_1589 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_6_), .Y(_11283_) );
	NAND2X1 NAND2X1_2072 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf7), .B(_11283_), .Y(_11284_) );
	NAND2X1 NAND2X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_11282_), .B(_11284_), .Y(_11285_) );
	NAND2X1 NAND2X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_11285_), .B(_11281_), .Y(_11286_) );
	NAND2X1 NAND2X1_2075 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_7_), .B(_11450__bF_buf3), .Y(_11287_) );
	NAND2X1 NAND2X1_2076 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(_11280_), .Y(_11288_) );
	NAND2X1 NAND2X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_11287_), .B(_11288_), .Y(_11289_) );
	NAND2X1 NAND2X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_11289_), .B(_11286_), .Y(_11290_) );
	OAI21X1 OAI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_11280_), .B(_11286_), .C(_11290_), .Y(divider_flipSign_rem_result_7_) );
	AOI22X1 AOI22X1_259 ( .gnd(gnd), .vdd(vdd), .A(_11461_), .B(_11468_), .C(_11473_), .D(_11474_), .Y(_11291_) );
	AOI22X1 AOI22X1_260 ( .gnd(gnd), .vdd(vdd), .A(_11282_), .B(_11284_), .C(_11287_), .D(_11288_), .Y(_11292_) );
	NAND2X1 NAND2X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_11291_), .B(_11292_), .Y(_11293_) );
	OAI21X1 OAI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_11466_), .B(_11293_), .C(divider_a_isNegative_bF_buf5), .Y(_11294_) );
	XNOR2X1 XNOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_11294_), .B(divider_flipSign_rem_operand_8_), .Y(divider_flipSign_rem_result_8_) );
	INVX1 INVX1_1590 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_9_), .Y(_11295_) );
	NOR2X1 NOR2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_11466_), .B(_11293_), .Y(_11296_) );
	NAND2X1 NAND2X1_2080 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_8_), .B(_11450__bF_buf2), .Y(_11297_) );
	INVX1 INVX1_1591 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_8_), .Y(_11298_) );
	NAND2X1 NAND2X1_2081 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(_11298_), .Y(_11299_) );
	NAND2X1 NAND2X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .B(_11299_), .Y(_11300_) );
	NAND2X1 NAND2X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_11300_), .B(_11296_), .Y(_11301_) );
	NAND2X1 NAND2X1_2084 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_9_), .B(_11450__bF_buf1), .Y(_11302_) );
	NAND2X1 NAND2X1_2085 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(_11295_), .Y(_11303_) );
	NAND2X1 NAND2X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_11302_), .B(_11303_), .Y(_11304_) );
	NAND2X1 NAND2X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_11304_), .B(_11301_), .Y(_11305_) );
	OAI21X1 OAI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_11295_), .B(_11301_), .C(_11305_), .Y(divider_flipSign_rem_result_9_) );
	OAI21X1 OAI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_9_), .B(_11301_), .C(divider_a_isNegative_bF_buf2), .Y(_11306_) );
	XNOR2X1 XNOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_11306_), .B(divider_flipSign_rem_operand_10_), .Y(divider_flipSign_rem_result_10_) );
	INVX1 INVX1_1592 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_11_), .Y(_11307_) );
	AOI22X1 AOI22X1_261 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .B(_11299_), .C(_11302_), .D(_11303_), .Y(_11308_) );
	NAND2X1 NAND2X1_2088 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_10_), .B(_11450__bF_buf0), .Y(_11309_) );
	INVX1 INVX1_1593 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_10_), .Y(_11310_) );
	NAND2X1 NAND2X1_2089 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(_11310_), .Y(_11311_) );
	NAND2X1 NAND2X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_11309_), .B(_11311_), .Y(_11312_) );
	NAND3X1 NAND3X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_11312_), .C(_11296_), .Y(_11313_) );
	NAND2X1 NAND2X1_2091 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_11_), .B(_11450__bF_buf4), .Y(_11314_) );
	NAND2X1 NAND2X1_2092 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(_11307_), .Y(_11315_) );
	NAND2X1 NAND2X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_11314_), .B(_11315_), .Y(_11316_) );
	NAND2X1 NAND2X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_11316_), .B(_11313_), .Y(_11317_) );
	OAI21X1 OAI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_11307_), .B(_11313_), .C(_11317_), .Y(divider_flipSign_rem_result_11_) );
	NAND2X1 NAND2X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_11296_), .Y(_11318_) );
	AOI22X1 AOI22X1_262 ( .gnd(gnd), .vdd(vdd), .A(_11309_), .B(_11311_), .C(_11314_), .D(_11315_), .Y(_11319_) );
	INVX1 INVX1_1594 ( .gnd(gnd), .vdd(vdd), .A(_11319_), .Y(_11320_) );
	OAI21X1 OAI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_11318_), .C(divider_a_isNegative_bF_buf8), .Y(_11321_) );
	XNOR2X1 XNOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_11321_), .B(divider_flipSign_rem_operand_12_), .Y(divider_flipSign_rem_result_12_) );
	INVX1 INVX1_1595 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_13_), .Y(_11322_) );
	NOR2X1 NOR2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_11318_), .Y(_11323_) );
	NAND2X1 NAND2X1_2096 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_12_), .B(_11450__bF_buf3), .Y(_11324_) );
	INVX1 INVX1_1596 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_12_), .Y(_11325_) );
	NAND2X1 NAND2X1_2097 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf7), .B(_11325_), .Y(_11326_) );
	NAND2X1 NAND2X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_11324_), .B(_11326_), .Y(_11327_) );
	NAND2X1 NAND2X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_11327_), .B(_11323_), .Y(_11328_) );
	NAND2X1 NAND2X1_2100 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_13_), .B(_11450__bF_buf2), .Y(_11329_) );
	NAND2X1 NAND2X1_2101 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(_11322_), .Y(_11330_) );
	NAND2X1 NAND2X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_11329_), .B(_11330_), .Y(_11331_) );
	NAND2X1 NAND2X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_11331_), .B(_11328_), .Y(_11332_) );
	OAI21X1 OAI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_11322_), .B(_11328_), .C(_11332_), .Y(divider_flipSign_rem_result_13_) );
	INVX1 INVX1_1597 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_14_), .Y(_11333_) );
	NAND3X1 NAND3X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_11319_), .C(_11296_), .Y(_11334_) );
	AOI22X1 AOI22X1_263 ( .gnd(gnd), .vdd(vdd), .A(_11324_), .B(_11326_), .C(_11329_), .D(_11330_), .Y(_11335_) );
	INVX1 INVX1_1598 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .Y(_11336_) );
	NOR2X1 NOR2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_11336_), .B(_11334_), .Y(_11337_) );
	NAND2X1 NAND2X1_2104 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_14_), .B(_11450__bF_buf1), .Y(_11338_) );
	NAND2X1 NAND2X1_2105 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(_11333_), .Y(_11339_) );
	NAND2X1 NAND2X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_11338_), .B(_11339_), .Y(_11340_) );
	AOI21X1 AOI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_11323_), .B(_11335_), .C(_11340_), .Y(_11341_) );
	AOI21X1 AOI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_11333_), .B(_11337_), .C(_11341_), .Y(divider_flipSign_rem_result_14_) );
	INVX1 INVX1_1599 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_15_), .Y(_11342_) );
	NAND2X1 NAND2X1_2107 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_15_), .B(_11450__bF_buf0), .Y(_11343_) );
	NAND2X1 NAND2X1_2108 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(_11342_), .Y(_11344_) );
	NAND2X1 NAND2X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_11343_), .B(_11344_), .Y(_11345_) );
	INVX1 INVX1_1600 ( .gnd(gnd), .vdd(vdd), .A(_11345_), .Y(_11346_) );
	NAND2X1 NAND2X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_11340_), .B(_11337_), .Y(_11347_) );
	MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_11346_), .B(_11342_), .S(_11347_), .Y(divider_flipSign_rem_result_15_) );
	NAND2X1 NAND2X1_2111 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_16_), .B(_11450__bF_buf4), .Y(_11348_) );
	NAND2X1 NAND2X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_11319_), .Y(_11349_) );
	AOI22X1 AOI22X1_264 ( .gnd(gnd), .vdd(vdd), .A(_11338_), .B(_11339_), .C(_11343_), .D(_11344_), .Y(_11350_) );
	NAND2X1 NAND2X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11350_), .Y(_11351_) );
	NOR2X1 NOR2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_11349_), .B(_11351_), .Y(_11352_) );
	AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_11352_), .B(_11296_), .Y(_11353_) );
	INVX1 INVX1_1601 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_16_), .Y(_11354_) );
	NAND2X1 NAND2X1_2114 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(_11354_), .Y(_11355_) );
	NAND2X1 NAND2X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_11348_), .B(_11355_), .Y(_11356_) );
	XNOR2X1 XNOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_11353_), .B(_11356_), .Y(_11357_) );
	OAI21X1 OAI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_11450__bF_buf3), .B(_11357_), .C(_11348_), .Y(divider_flipSign_rem_result_16_) );
	INVX1 INVX1_1602 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_17_), .Y(_11358_) );
	NAND2X1 NAND2X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_11308_), .B(_11350_), .Y(_11359_) );
	NAND2X1 NAND2X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_11319_), .B(_11335_), .Y(_11360_) );
	NOR2X1 NOR2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_11359_), .B(_11360_), .Y(_11361_) );
	AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_11361_), .B(_11296_), .Y(_11362_) );
	NAND2X1 NAND2X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_11356_), .B(_11362_), .Y(_11363_) );
	INVX1 INVX1_1603 ( .gnd(gnd), .vdd(vdd), .A(_11353_), .Y(_11364_) );
	INVX1 INVX1_1604 ( .gnd(gnd), .vdd(vdd), .A(_11356_), .Y(_11365_) );
	NAND2X1 NAND2X1_2119 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_17_), .B(_11450__bF_buf2), .Y(_11366_) );
	NAND2X1 NAND2X1_2120 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(_11358_), .Y(_11367_) );
	NAND2X1 NAND2X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_11366_), .B(_11367_), .Y(_11368_) );
	OAI21X1 OAI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_11365_), .B(_11364_), .C(_11368_), .Y(_11369_) );
	OAI21X1 OAI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_11358_), .B(_11363_), .C(_11369_), .Y(divider_flipSign_rem_result_17_) );
	INVX1 INVX1_1605 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_18_), .Y(_11370_) );
	AOI22X1 AOI22X1_265 ( .gnd(gnd), .vdd(vdd), .A(_11348_), .B(_11355_), .C(_11366_), .D(_11367_), .Y(_11371_) );
	AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_11362_), .B(_11371_), .Y(_11372_) );
	NAND2X1 NAND2X1_2122 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_18_), .B(_11450__bF_buf1), .Y(_11373_) );
	NAND2X1 NAND2X1_2123 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(_11370_), .Y(_11374_) );
	NAND2X1 NAND2X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_11373_), .B(_11374_), .Y(_11375_) );
	NOR2X1 NOR2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_11375_), .B(_11372_), .Y(_11376_) );
	AOI21X1 AOI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_11370_), .B(_11372_), .C(_11376_), .Y(divider_flipSign_rem_result_18_) );
	INVX1 INVX1_1606 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_19_), .Y(_11377_) );
	NAND2X1 NAND2X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_11375_), .B(_11372_), .Y(_11378_) );
	XOR2X1 XOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(divider_flipSign_rem_operand_19_), .Y(_11379_) );
	NAND2X1 NAND2X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_11379_), .B(_11378_), .Y(_11380_) );
	OAI21X1 OAI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_11377_), .B(_11378_), .C(_11380_), .Y(divider_flipSign_rem_result_19_) );
	NAND3X1 NAND3X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_11375_), .B(_11379_), .C(_11371_), .Y(_11381_) );
	OAI21X1 OAI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .B(_11364_), .C(divider_a_isNegative_bF_buf8), .Y(_11382_) );
	XNOR2X1 XNOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_11382_), .B(divider_flipSign_rem_operand_20_), .Y(divider_flipSign_rem_result_20_) );
	INVX1 INVX1_1607 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_21_), .Y(_11383_) );
	NAND2X1 NAND2X1_2127 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_21_), .B(_11450__bF_buf0), .Y(_11384_) );
	NAND2X1 NAND2X1_2128 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf7), .B(_11383_), .Y(_11385_) );
	AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_11384_), .B(_11385_), .Y(_11386_) );
	INVX1 INVX1_1608 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .Y(_11387_) );
	NAND2X1 NAND2X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_11387_), .B(_11362_), .Y(_11388_) );
	NAND2X1 NAND2X1_2130 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_20_), .B(_11450__bF_buf4), .Y(_11389_) );
	INVX1 INVX1_1609 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_20_), .Y(_11390_) );
	NAND2X1 NAND2X1_2131 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(_11390_), .Y(_11391_) );
	AOI21X1 AOI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_11389_), .B(_11391_), .C(_11388_), .Y(_11392_) );
	MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_11383_), .B(_11386_), .S(_11392_), .Y(divider_flipSign_rem_result_21_) );
	INVX1 INVX1_1610 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_22_), .Y(_11393_) );
	NAND2X1 NAND2X1_2132 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_22_), .B(_11450__bF_buf3), .Y(_11394_) );
	NAND2X1 NAND2X1_2133 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(_11393_), .Y(_11395_) );
	NAND2X1 NAND2X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_11394_), .B(_11395_), .Y(_11396_) );
	INVX1 INVX1_1611 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .Y(_11397_) );
	AOI22X1 AOI22X1_266 ( .gnd(gnd), .vdd(vdd), .A(_11389_), .B(_11391_), .C(_11384_), .D(_11385_), .Y(_11398_) );
	INVX1 INVX1_1612 ( .gnd(gnd), .vdd(vdd), .A(_11398_), .Y(_11399_) );
	NOR2X1 NOR2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_11399_), .B(_11388_), .Y(_11400_) );
	MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11397_), .S(_11400_), .Y(divider_flipSign_rem_result_22_) );
	XOR2X1 XOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(divider_flipSign_rem_operand_23_), .Y(_11401_) );
	INVX1 INVX1_1613 ( .gnd(gnd), .vdd(vdd), .A(_11401_), .Y(_11402_) );
	NAND2X1 NAND2X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_11387_), .B(_11353_), .Y(_11403_) );
	NOR3X1 NOR3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_11397_), .B(_11399_), .C(_11403_), .Y(_11404_) );
	NAND3X1 NAND3X1_2306 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_23_), .B(_11396_), .C(_11400_), .Y(_11405_) );
	OAI21X1 OAI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_11402_), .B(_11404_), .C(_11405_), .Y(divider_flipSign_rem_result_23_) );
	NAND2X1 NAND2X1_2136 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_24_), .B(_11450__bF_buf2), .Y(_11406_) );
	INVX1 INVX1_1614 ( .gnd(gnd), .vdd(vdd), .A(_11406_), .Y(_11407_) );
	NOR2X1 NOR2X1_745 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_24_), .B(_11450__bF_buf1), .Y(_11408_) );
	OR2X2 OR2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_11407_), .B(_11408_), .Y(_11409_) );
	NAND3X1 NAND3X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11401_), .C(_11398_), .Y(_11410_) );
	NOR2X1 NOR2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_11381_), .B(_11410_), .Y(_11411_) );
	NAND3X1 NAND3X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_11296_), .B(_11352_), .C(_11411_), .Y(_11412_) );
	XOR2X1 XOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_11412_), .B(_11409_), .Y(_11413_) );
	OAI21X1 OAI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_11450__bF_buf0), .B(_11413_), .C(_11406_), .Y(divider_flipSign_rem_result_24_) );
	OAI21X1 OAI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_24_), .B(_11412_), .C(divider_a_isNegative_bF_buf3), .Y(_11414_) );
	XNOR2X1 XNOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_11414_), .B(divider_flipSign_rem_operand_25_), .Y(divider_flipSign_rem_result_25_) );
	XOR2X1 XOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf2), .B(divider_flipSign_rem_operand_25_), .Y(_11415_) );
	OAI21X1 OAI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_11408_), .B(_11407_), .C(_11415_), .Y(_11416_) );
	OAI21X1 OAI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_11416_), .B(_11412_), .C(divider_a_isNegative_bF_buf1), .Y(_11417_) );
	XNOR2X1 XNOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_11417_), .B(divider_flipSign_rem_operand_26_), .Y(divider_flipSign_rem_result_26_) );
	XOR2X1 XOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf0), .B(divider_flipSign_rem_operand_27_), .Y(_11418_) );
	INVX1 INVX1_1615 ( .gnd(gnd), .vdd(vdd), .A(_11418_), .Y(_11419_) );
	NOR2X1 NOR2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_11416_), .B(_11412_), .Y(_11420_) );
	XOR2X1 XOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf8), .B(divider_flipSign_rem_operand_26_), .Y(_11421_) );
	NAND2X1 NAND2X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_11421_), .B(_11420_), .Y(_11422_) );
	NOR2X1 NOR2X1_748 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_27_), .B(_11422_), .Y(_11423_) );
	AOI21X1 AOI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_11419_), .B(_11422_), .C(_11423_), .Y(divider_flipSign_rem_result_27_) );
	INVX1 INVX1_1616 ( .gnd(gnd), .vdd(vdd), .A(_11416_), .Y(_11424_) );
	AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_11421_), .B(_11418_), .Y(_11425_) );
	NAND2X1 NAND2X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_11425_), .B(_11424_), .Y(_11426_) );
	OAI21X1 OAI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_11426_), .B(_11412_), .C(divider_a_isNegative_bF_buf7), .Y(_11427_) );
	XNOR2X1 XNOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_11427_), .B(divider_flipSign_rem_operand_28_), .Y(divider_flipSign_rem_result_28_) );
	XOR2X1 XOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf6), .B(divider_flipSign_rem_operand_29_), .Y(_11428_) );
	INVX1 INVX1_1617 ( .gnd(gnd), .vdd(vdd), .A(_11428_), .Y(_11429_) );
	NOR2X1 NOR2X1_749 ( .gnd(gnd), .vdd(vdd), .A(_11426_), .B(_11412_), .Y(_11430_) );
	XNOR2X1 XNOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf5), .B(divider_flipSign_rem_operand_28_), .Y(_11431_) );
	INVX1 INVX1_1618 ( .gnd(gnd), .vdd(vdd), .A(_11431_), .Y(_11432_) );
	NAND2X1 NAND2X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_11432_), .B(_11430_), .Y(_11433_) );
	NOR2X1 NOR2X1_750 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_29_), .B(_11433_), .Y(_11434_) );
	AOI21X1 AOI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11433_), .C(_11434_), .Y(divider_flipSign_rem_result_29_) );
	INVX1 INVX1_1619 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_30_), .Y(_11435_) );
	NAND2X1 NAND2X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_11428_), .B(_11432_), .Y(_11436_) );
	NOR3X1 NOR3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_11426_), .B(_11436_), .C(_11412_), .Y(_11437_) );
	OAI21X1 OAI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_11450__bF_buf4), .B(_11437_), .C(_11435_), .Y(_11438_) );
	INVX1 INVX1_1620 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .Y(_11439_) );
	NAND2X1 NAND2X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_11439_), .B(_11430_), .Y(_11440_) );
	NAND3X1 NAND3X1_2309 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf4), .B(divider_flipSign_rem_operand_30_), .C(_11440_), .Y(_11441_) );
	AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_11441_), .B(_11438_), .Y(divider_flipSign_rem_result_30_) );
	INVX1 INVX1_1621 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_31_), .Y(_11442_) );
	NAND3X1 NAND3X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_11435_), .B(_11439_), .C(_11430_), .Y(_11443_) );
	NAND3X1 NAND3X1_2311 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf3), .B(_11442_), .C(_11443_), .Y(_11444_) );
	INVX1 INVX1_1622 ( .gnd(gnd), .vdd(vdd), .A(_11426_), .Y(_11445_) );
	NAND3X1 NAND3X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_11411_), .B(_11445_), .C(_11353_), .Y(_11446_) );
	OAI21X1 OAI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .B(_11446_), .C(divider_a_isNegative_bF_buf2), .Y(_11447_) );
	NAND2X1 NAND2X1_2142 ( .gnd(gnd), .vdd(vdd), .A(divider_a_isNegative_bF_buf1), .B(divider_flipSign_rem_operand_30_), .Y(_11448_) );
	NAND3X1 NAND3X1_2313 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_31_), .B(_11448_), .C(_11447_), .Y(_11449_) );
	NAND2X1 NAND2X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_11444_), .B(_11449_), .Y(divider_flipSign_rem_result_31_) );
	BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(divider_flipSign_rem_operand_0_), .Y(divider_flipSign_rem_result_0_) );
	OR2X2 OR2X2_126 ( .gnd(gnd), .vdd(vdd), .A(frameWriteController_writebackState), .B(executeState), .Y(frameWriteController_result_we) );
	INVX1 INVX1_1623 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[14]), .Y(_11478_) );
	NOR2X1 NOR2X1_751 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[3]), .B(instructionIn[2]), .Y(_11479_) );
	AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[1]), .B(instructionIn[0]), .Y(_11480_) );
	NAND2X1 NAND2X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_11479_), .B(_11480_), .Y(_11481_) );
	INVX1 INVX1_1624 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[6]), .Y(_11482_) );
	NAND3X1 NAND3X1_2314 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[5]), .B(instructionIn[4]), .C(_11482_), .Y(_11483_) );
	NOR2X1 NOR2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_11483_), .B(_11481_), .Y(_11484_) );
	NOR2X1 NOR2X1_753 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[13]), .B(instructionIn[12]), .Y(_11485_) );
	NAND3X1 NAND3X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_11478_), .B(_11485_), .C(_11484_), .Y(_11486_) );
	NOR2X1 NOR2X1_754 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[28]), .B(instructionIn[27]), .Y(_11487_) );
	NOR2X1 NOR2X1_755 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[25]), .B(instructionIn[26]), .Y(_11488_) );
	INVX1 INVX1_1625 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[30]), .Y(_11489_) );
	INVX1 INVX1_1626 ( .gnd(gnd), .vdd(vdd), .A(instructionIn_31_bF_buf3), .Y(_11490_) );
	INVX1 INVX1_1627 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[29]), .Y(_11491_) );
	NAND2X1 NAND2X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_11490_), .B(_11491_), .Y(_11492_) );
	NOR2X1 NOR2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_11489_), .B(_11492_), .Y(_11493_) );
	NAND3X1 NAND3X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_11487_), .B(_11488_), .C(_11493_), .Y(_11494_) );
	NOR2X1 NOR2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_11494_), .B(_11486_), .Y(instructionDecoder_sub_flag) );
	NOR2X1 NOR2X1_758 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[6]), .B(instructionIn[5]), .Y(_11495_) );
	NAND2X1 NAND2X1_2146 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[4]), .B(_11495_), .Y(_11496_) );
	NOR2X1 NOR2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_11496_), .B(_11481_), .Y(_11497_) );
	INVX1 INVX1_1628 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[13]), .Y(_11498_) );
	AOI21X1 AOI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_11498_), .B(instructionIn[12]), .C(instructionIn[14]), .Y(_11499_) );
	AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11499_), .Y(immediateSelect_decodeOut) );
	INVX1 INVX1_1629 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[12]), .Y(_11500_) );
	NAND3X1 NAND3X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_11489_), .B(_11490_), .C(_11491_), .Y(_11501_) );
	INVX1 INVX1_1630 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[26]), .Y(_11502_) );
	NAND3X1 NAND3X1_2318 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[25]), .B(_11502_), .C(_11487_), .Y(_11503_) );
	NOR2X1 NOR2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_11501_), .B(_11503_), .Y(_11504_) );
	NAND3X1 NAND3X1_2319 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[14]), .B(_11484_), .C(_11504_), .Y(_11505_) );
	NAND3X1 NAND3X1_2320 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[13]), .B(instructionIn[12]), .C(_11478_), .Y(_11506_) );
	INVX1 INVX1_1631 ( .gnd(gnd), .vdd(vdd), .A(_11506_), .Y(_11507_) );
	NAND2X1 NAND2X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_11487_), .B(_11488_), .Y(_11508_) );
	NOR2X1 NOR2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_11501_), .B(_11508_), .Y(_11509_) );
	NOR3X1 NOR3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_11483_), .B(_11506_), .C(_11481_), .Y(_11510_) );
	AOI22X1 AOI22X1_267 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11507_), .C(_11509_), .D(_11510_), .Y(_11511_) );
	OAI21X1 OAI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_11500_), .B(_11505_), .C(_11511_), .Y(instructionDecoder_unsignedSelect) );
	INVX1 INVX1_1632 ( .gnd(gnd), .vdd(vdd), .A(_11504_), .Y(_11512_) );
	OAI22X1 OAI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_11486_), .B(_11512_), .C(_11498_), .D(_11505_), .Y(instructionDecoder_resultSelect_0_) );
	NAND2X1 NAND2X1_2148 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[13]), .B(_11478_), .Y(_11513_) );
	INVX1 INVX1_1633 ( .gnd(gnd), .vdd(vdd), .A(_11513_), .Y(_11514_) );
	AOI22X1 AOI22X1_268 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11514_), .C(_11509_), .D(_11510_), .Y(_11515_) );
	NOR2X1 NOR2X1_762 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[12]), .B(_11513_), .Y(_11516_) );
	NAND3X1 NAND3X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_11516_), .B(_11509_), .C(_11484_), .Y(_11517_) );
	NAND3X1 NAND3X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_11505_), .B(_11517_), .C(_11515_), .Y(instructionDecoder_resultSelect_1_) );
	NAND2X1 NAND2X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_11517_), .B(_11515_), .Y(instructionDecoder_resultSelect_2_) );
	NAND2X1 NAND2X1_2150 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(aLoc_we), .Y(_11529_) );
	INVX1 INVX1_1634 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11530_) );
	NAND2X1 NAND2X1_2151 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeEnable_out), .B(_11530_), .Y(_11531_) );
	AOI21X1 AOI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_11531_), .B(_11529_), .C(reset_bF_buf10), .Y(_11527_) );
	NAND2X1 NAND2X1_2152 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[7]), .B(aLoc_we), .Y(_11532_) );
	INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11533_) );
	NAND2X1 NAND2X1_2153 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_0_), .B(_11533_), .Y(_11534_) );
	AOI21X1 AOI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_11534_), .B(_11532_), .C(reset_bF_buf9), .Y(_11528__0_) );
	NAND2X1 NAND2X1_2154 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[8]), .Y(_11535_) );
	NAND2X1 NAND2X1_2155 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_1_), .B(_11533_), .Y(_11536_) );
	AOI21X1 AOI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .B(_11535_), .C(reset_bF_buf8), .Y(_11528__1_) );
	NAND2X1 NAND2X1_2156 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[9]), .Y(_11537_) );
	NAND2X1 NAND2X1_2157 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_2_), .B(_11533_), .Y(_11538_) );
	AOI21X1 AOI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_11538_), .B(_11537_), .C(reset_bF_buf7), .Y(_11528__2_) );
	NAND2X1 NAND2X1_2158 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[10]), .Y(_11539_) );
	NAND2X1 NAND2X1_2159 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_3_), .B(_11533_), .Y(_11540_) );
	AOI21X1 AOI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_11540_), .B(_11539_), .C(reset_bF_buf6), .Y(_11528__3_) );
	NAND2X1 NAND2X1_2160 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[11]), .Y(_11541_) );
	NAND2X1 NAND2X1_2161 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_4_), .B(_11533_), .Y(_11542_) );
	AOI21X1 AOI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_11542_), .B(_11541_), .C(reset_bF_buf5), .Y(_11528__4_) );
	NAND2X1 NAND2X1_2162 ( .gnd(gnd), .vdd(vdd), .A(instructionDecoder_resultSelect_0_), .B(aLoc_we), .Y(_11543_) );
	INVX1 INVX1_1635 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11544_) );
	NAND2X1 NAND2X1_2163 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_0_), .B(_11544_), .Y(_11545_) );
	AOI21X1 AOI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_11545_), .B(_11543_), .C(reset_bF_buf4), .Y(_11524__0_) );
	NAND2X1 NAND2X1_2164 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionDecoder_resultSelect_1_), .Y(_11546_) );
	NAND2X1 NAND2X1_2165 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_1_), .B(_11544_), .Y(_11547_) );
	AOI21X1 AOI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_11547_), .B(_11546_), .C(reset_bF_buf3), .Y(_11524__1_) );
	NAND2X1 NAND2X1_2166 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionDecoder_resultSelect_2_), .Y(_11548_) );
	NAND2X1 NAND2X1_2167 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_resultSelect_out_2_), .B(_11544_), .Y(_11549_) );
	AOI21X1 AOI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_11549_), .B(_11548_), .C(reset_bF_buf2), .Y(_11524__2_) );
	NAND2X1 NAND2X1_2168 ( .gnd(gnd), .vdd(vdd), .A(instructionDecoder_sub_flag), .B(aLoc_we), .Y(_11550_) );
	INVX1 INVX1_1636 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11551_) );
	NAND2X1 NAND2X1_2169 ( .gnd(gnd), .vdd(vdd), .A(adder_subtract_bF_buf2), .B(_11551_), .Y(_11552_) );
	AOI21X1 AOI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_11552_), .B(_11550_), .C(reset_bF_buf1), .Y(_11525_) );
	NAND2X1 NAND2X1_2170 ( .gnd(gnd), .vdd(vdd), .A(instructionDecoder_unsignedSelect), .B(aLoc_we), .Y(_11553_) );
	INVX1 INVX1_1637 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11554_) );
	NAND2X1 NAND2X1_2171 ( .gnd(gnd), .vdd(vdd), .A(comparator_unsignedEn), .B(_11554_), .Y(_11555_) );
	AOI21X1 AOI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_11555_), .B(_11553_), .C(reset_bF_buf0), .Y(_11526_) );
	NAND2X1 NAND2X1_2172 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_decodeOut), .B(aLoc_we), .Y(_11556_) );
	INVX1 INVX1_1638 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11557_) );
	NAND2X1 NAND2X1_2173 ( .gnd(gnd), .vdd(vdd), .A(immediateSelect_frameOut_bF_buf7), .B(_11557_), .Y(_11558_) );
	AOI21X1 AOI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_11558_), .B(_11556_), .C(reset_bF_buf10), .Y(_11522_) );
	NAND2X1 NAND2X1_2174 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[20]), .B(aLoc_we), .Y(_11559_) );
	INVX8 INVX8_45 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11560_) );
	NAND2X1 NAND2X1_2175 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_0_), .B(_11560__bF_buf4), .Y(_11561_) );
	AOI21X1 AOI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_11561_), .B(_11559_), .C(reset_bF_buf9), .Y(_11523__0_) );
	NAND2X1 NAND2X1_2176 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[21]), .Y(_11562_) );
	NAND2X1 NAND2X1_2177 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_1_), .B(_11560__bF_buf3), .Y(_11563_) );
	AOI21X1 AOI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_11563_), .B(_11562_), .C(reset_bF_buf8), .Y(_11523__1_) );
	NAND2X1 NAND2X1_2178 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[22]), .Y(_11564_) );
	NAND2X1 NAND2X1_2179 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_2_), .B(_11560__bF_buf2), .Y(_11565_) );
	AOI21X1 AOI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_11565_), .B(_11564_), .C(reset_bF_buf7), .Y(_11523__2_) );
	NAND2X1 NAND2X1_2180 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[23]), .Y(_11566_) );
	NAND2X1 NAND2X1_2181 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_3_), .B(_11560__bF_buf1), .Y(_11567_) );
	AOI21X1 AOI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_11567_), .B(_11566_), .C(reset_bF_buf6), .Y(_11523__3_) );
	NAND2X1 NAND2X1_2182 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[24]), .Y(_11568_) );
	NAND2X1 NAND2X1_2183 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_4_), .B(_11560__bF_buf0), .Y(_11569_) );
	AOI21X1 AOI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_11569_), .B(_11568_), .C(reset_bF_buf5), .Y(_11523__4_) );
	NAND2X1 NAND2X1_2184 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[25]), .Y(_11570_) );
	NAND2X1 NAND2X1_2185 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_5_), .B(_11560__bF_buf4), .Y(_11571_) );
	AOI21X1 AOI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_11571_), .B(_11570_), .C(reset_bF_buf4), .Y(_11523__5_) );
	NAND2X1 NAND2X1_2186 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[26]), .Y(_11572_) );
	NAND2X1 NAND2X1_2187 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_6_), .B(_11560__bF_buf3), .Y(_11573_) );
	AOI21X1 AOI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_11573_), .B(_11572_), .C(reset_bF_buf3), .Y(_11523__6_) );
	NAND2X1 NAND2X1_2188 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[27]), .Y(_11574_) );
	NAND2X1 NAND2X1_2189 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_7_), .B(_11560__bF_buf2), .Y(_11575_) );
	AOI21X1 AOI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_11575_), .B(_11574_), .C(reset_bF_buf2), .Y(_11523__7_) );
	NAND2X1 NAND2X1_2190 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[28]), .Y(_11576_) );
	NAND2X1 NAND2X1_2191 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_8_), .B(_11560__bF_buf1), .Y(_11577_) );
	AOI21X1 AOI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_11577_), .B(_11576_), .C(reset_bF_buf1), .Y(_11523__8_) );
	NAND2X1 NAND2X1_2192 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[29]), .Y(_11578_) );
	NAND2X1 NAND2X1_2193 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_9_), .B(_11560__bF_buf0), .Y(_11579_) );
	AOI21X1 AOI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_11579_), .B(_11578_), .C(reset_bF_buf0), .Y(_11523__9_) );
	NAND2X1 NAND2X1_2194 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[30]), .Y(_11580_) );
	NAND2X1 NAND2X1_2195 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_10_), .B(_11560__bF_buf4), .Y(_11581_) );
	AOI21X1 AOI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_11581_), .B(_11580_), .C(reset_bF_buf10), .Y(_11523__10_) );
	NAND2X1 NAND2X1_2196 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf2), .Y(_11582_) );
	NAND2X1 NAND2X1_2197 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_11_), .B(_11560__bF_buf3), .Y(_11583_) );
	AOI21X1 AOI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_11583_), .B(_11582_), .C(reset_bF_buf9), .Y(_11523__11_) );
	NAND2X1 NAND2X1_2198 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf1), .Y(_11584_) );
	NAND2X1 NAND2X1_2199 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_12_), .B(_11560__bF_buf2), .Y(_11585_) );
	AOI21X1 AOI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_11585_), .B(_11584_), .C(reset_bF_buf8), .Y(_11523__12_) );
	NAND2X1 NAND2X1_2200 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf0), .Y(_11586_) );
	NAND2X1 NAND2X1_2201 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_13_), .B(_11560__bF_buf1), .Y(_11587_) );
	AOI21X1 AOI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_11587_), .B(_11586_), .C(reset_bF_buf7), .Y(_11523__13_) );
	NAND2X1 NAND2X1_2202 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf3), .Y(_11588_) );
	NAND2X1 NAND2X1_2203 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_14_), .B(_11560__bF_buf0), .Y(_11589_) );
	AOI21X1 AOI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_11589_), .B(_11588_), .C(reset_bF_buf6), .Y(_11523__14_) );
	NAND2X1 NAND2X1_2204 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf2), .Y(_11590_) );
	NAND2X1 NAND2X1_2205 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_15_), .B(_11560__bF_buf4), .Y(_11591_) );
	AOI21X1 AOI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_11591_), .B(_11590_), .C(reset_bF_buf5), .Y(_11523__15_) );
	NAND2X1 NAND2X1_2206 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf1), .Y(_11592_) );
	NAND2X1 NAND2X1_2207 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_16_), .B(_11560__bF_buf3), .Y(_11593_) );
	AOI21X1 AOI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_11593_), .B(_11592_), .C(reset_bF_buf4), .Y(_11523__16_) );
	NAND2X1 NAND2X1_2208 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf0), .Y(_11594_) );
	NAND2X1 NAND2X1_2209 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_17_), .B(_11560__bF_buf2), .Y(_11595_) );
	AOI21X1 AOI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_11595_), .B(_11594_), .C(reset_bF_buf3), .Y(_11523__17_) );
	NAND2X1 NAND2X1_2210 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf3), .Y(_11596_) );
	NAND2X1 NAND2X1_2211 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_18_), .B(_11560__bF_buf1), .Y(_11597_) );
	AOI21X1 AOI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_11597_), .B(_11596_), .C(reset_bF_buf2), .Y(_11523__18_) );
	NAND2X1 NAND2X1_2212 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf2), .Y(_11598_) );
	NAND2X1 NAND2X1_2213 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_19_), .B(_11560__bF_buf0), .Y(_11599_) );
	AOI21X1 AOI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_11599_), .B(_11598_), .C(reset_bF_buf1), .Y(_11523__19_) );
	NAND2X1 NAND2X1_2214 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf1), .Y(_11600_) );
	NAND2X1 NAND2X1_2215 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_20_), .B(_11560__bF_buf4), .Y(_11601_) );
	AOI21X1 AOI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_11601_), .B(_11600_), .C(reset_bF_buf0), .Y(_11523__20_) );
	NAND2X1 NAND2X1_2216 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf0), .Y(_11602_) );
	NAND2X1 NAND2X1_2217 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_21_), .B(_11560__bF_buf3), .Y(_11603_) );
	AOI21X1 AOI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_11603_), .B(_11602_), .C(reset_bF_buf10), .Y(_11523__21_) );
	NAND2X1 NAND2X1_2218 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf3), .Y(_11604_) );
	NAND2X1 NAND2X1_2219 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_22_), .B(_11560__bF_buf2), .Y(_11605_) );
	AOI21X1 AOI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_11605_), .B(_11604_), .C(reset_bF_buf9), .Y(_11523__22_) );
	NAND2X1 NAND2X1_2220 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf2), .Y(_11606_) );
	NAND2X1 NAND2X1_2221 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_23_), .B(_11560__bF_buf1), .Y(_11607_) );
	AOI21X1 AOI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_11606_), .C(reset_bF_buf8), .Y(_11523__23_) );
	NAND2X1 NAND2X1_2222 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf1), .Y(_11608_) );
	NAND2X1 NAND2X1_2223 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_24_), .B(_11560__bF_buf0), .Y(_11609_) );
	AOI21X1 AOI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_11609_), .B(_11608_), .C(reset_bF_buf7), .Y(_11523__24_) );
	NAND2X1 NAND2X1_2224 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf0), .Y(_11610_) );
	NAND2X1 NAND2X1_2225 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_25_), .B(_11560__bF_buf4), .Y(_11611_) );
	AOI21X1 AOI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_11611_), .B(_11610_), .C(reset_bF_buf6), .Y(_11523__25_) );
	NAND2X1 NAND2X1_2226 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf3), .Y(_11612_) );
	NAND2X1 NAND2X1_2227 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_26_), .B(_11560__bF_buf3), .Y(_11613_) );
	AOI21X1 AOI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_11613_), .B(_11612_), .C(reset_bF_buf5), .Y(_11523__26_) );
	NAND2X1 NAND2X1_2228 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf2), .Y(_11614_) );
	NAND2X1 NAND2X1_2229 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_27_), .B(_11560__bF_buf2), .Y(_11615_) );
	AOI21X1 AOI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_11615_), .B(_11614_), .C(reset_bF_buf4), .Y(_11523__27_) );
	NAND2X1 NAND2X1_2230 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf1), .Y(_11616_) );
	NAND2X1 NAND2X1_2231 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_28_), .B(_11560__bF_buf1), .Y(_11617_) );
	AOI21X1 AOI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_11617_), .B(_11616_), .C(reset_bF_buf3), .Y(_11523__28_) );
	NAND2X1 NAND2X1_2232 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf0), .Y(_11618_) );
	NAND2X1 NAND2X1_2233 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_29_), .B(_11560__bF_buf0), .Y(_11619_) );
	AOI21X1 AOI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_11619_), .B(_11618_), .C(reset_bF_buf2), .Y(_11523__29_) );
	NAND2X1 NAND2X1_2234 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf3), .Y(_11620_) );
	NAND2X1 NAND2X1_2235 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_30_), .B(_11560__bF_buf4), .Y(_11621_) );
	AOI21X1 AOI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_11621_), .B(_11620_), .C(reset_bF_buf1), .Y(_11523__30_) );
	NAND2X1 NAND2X1_2236 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn_31_bF_buf2), .Y(_11622_) );
	NAND2X1 NAND2X1_2237 ( .gnd(gnd), .vdd(vdd), .A(immediateVal_frameOut_31_), .B(_11560__bF_buf3), .Y(_11623_) );
	AOI21X1 AOI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_11623_), .B(_11622_), .C(reset_bF_buf0), .Y(_11523__31_) );
	NAND2X1 NAND2X1_2238 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[20]), .B(aLoc_we), .Y(_11624_) );
	INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11625_) );
	NAND2X1 NAND2X1_2239 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_0_), .B(_11625_), .Y(_11626_) );
	AOI21X1 AOI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_11626_), .B(_11624_), .C(reset_bF_buf10), .Y(_11520__0_) );
	NAND2X1 NAND2X1_2240 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[21]), .Y(_11627_) );
	NAND2X1 NAND2X1_2241 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .B(_11625_), .Y(_11628_) );
	AOI21X1 AOI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_11628_), .B(_11627_), .C(reset_bF_buf9), .Y(_11520__1_) );
	NAND2X1 NAND2X1_2242 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[22]), .Y(_11629_) );
	NAND2X1 NAND2X1_2243 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_2_), .B(_11625_), .Y(_11630_) );
	AOI21X1 AOI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_11630_), .B(_11629_), .C(reset_bF_buf8), .Y(_11520__2_) );
	NAND2X1 NAND2X1_2244 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[23]), .Y(_11631_) );
	NAND2X1 NAND2X1_2245 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_3_), .B(_11625_), .Y(_11632_) );
	AOI21X1 AOI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_11632_), .B(_11631_), .C(reset_bF_buf7), .Y(_11520__3_) );
	NAND2X1 NAND2X1_2246 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[24]), .Y(_11633_) );
	NAND2X1 NAND2X1_2247 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf6), .B(_11625_), .Y(_11634_) );
	AOI21X1 AOI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_11634_), .B(_11633_), .C(reset_bF_buf6), .Y(_11520__4_) );
	NAND2X1 NAND2X1_2248 ( .gnd(gnd), .vdd(vdd), .A(bOperand_frameIn_0_), .B(aOperand_we), .Y(_11635_) );
	INVX8 INVX8_46 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .Y(_11636_) );
	NAND2X1 NAND2X1_2249 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(_11636__bF_buf4), .Y(_11637_) );
	AOI21X1 AOI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_11637_), .B(_11635_), .C(reset_bF_buf5), .Y(_11521__0_) );
	NAND2X1 NAND2X1_2250 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_1_), .Y(_11638_) );
	NAND2X1 NAND2X1_2251 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(_11636__bF_buf3), .Y(_11639_) );
	AOI21X1 AOI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_11639_), .B(_11638_), .C(reset_bF_buf4), .Y(_11521__1_) );
	NAND2X1 NAND2X1_2252 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_2_), .Y(_11640_) );
	NAND2X1 NAND2X1_2253 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf1), .B(_11636__bF_buf2), .Y(_11641_) );
	AOI21X1 AOI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_11641_), .B(_11640_), .C(reset_bF_buf3), .Y(_11521__2_) );
	NAND2X1 NAND2X1_2254 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_3_), .Y(_11642_) );
	NAND2X1 NAND2X1_2255 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf3), .B(_11636__bF_buf1), .Y(_11643_) );
	AOI21X1 AOI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_11643_), .B(_11642_), .C(reset_bF_buf2), .Y(_11521__3_) );
	NAND2X1 NAND2X1_2256 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_4_), .Y(_11644_) );
	NAND2X1 NAND2X1_2257 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .B(_11636__bF_buf0), .Y(_11645_) );
	AOI21X1 AOI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_11645_), .B(_11644_), .C(reset_bF_buf1), .Y(_11521__4_) );
	NAND2X1 NAND2X1_2258 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_5_), .Y(_11646_) );
	NAND2X1 NAND2X1_2259 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf1), .B(_11636__bF_buf4), .Y(_11647_) );
	AOI21X1 AOI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_11647_), .B(_11646_), .C(reset_bF_buf0), .Y(_11521__5_) );
	NAND2X1 NAND2X1_2260 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_6_), .Y(_11648_) );
	NAND2X1 NAND2X1_2261 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf3), .B(_11636__bF_buf3), .Y(_11649_) );
	AOI21X1 AOI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_11649_), .B(_11648_), .C(reset_bF_buf10), .Y(_11521__6_) );
	NAND2X1 NAND2X1_2262 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_7_), .Y(_11650_) );
	NAND2X1 NAND2X1_2263 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf4), .B(_11636__bF_buf2), .Y(_11651_) );
	AOI21X1 AOI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_11651_), .B(_11650_), .C(reset_bF_buf9), .Y(_11521__7_) );
	NAND2X1 NAND2X1_2264 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_8_), .Y(_11652_) );
	NAND2X1 NAND2X1_2265 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf1), .B(_11636__bF_buf1), .Y(_11653_) );
	AOI21X1 AOI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_11653_), .B(_11652_), .C(reset_bF_buf8), .Y(_11521__8_) );
	NAND2X1 NAND2X1_2266 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_9_), .Y(_11654_) );
	NAND2X1 NAND2X1_2267 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf2), .B(_11636__bF_buf0), .Y(_11655_) );
	AOI21X1 AOI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_11655_), .B(_11654_), .C(reset_bF_buf7), .Y(_11521__9_) );
	NAND2X1 NAND2X1_2268 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_10_), .Y(_11656_) );
	NAND2X1 NAND2X1_2269 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf0), .B(_11636__bF_buf4), .Y(_11657_) );
	AOI21X1 AOI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_11657_), .B(_11656_), .C(reset_bF_buf6), .Y(_11521__10_) );
	NAND2X1 NAND2X1_2270 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_11_), .Y(_11658_) );
	NAND2X1 NAND2X1_2271 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf0), .B(_11636__bF_buf3), .Y(_11659_) );
	AOI21X1 AOI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_11659_), .B(_11658_), .C(reset_bF_buf5), .Y(_11521__11_) );
	NAND2X1 NAND2X1_2272 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_12_), .Y(_11660_) );
	NAND2X1 NAND2X1_2273 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf3), .B(_11636__bF_buf2), .Y(_11661_) );
	AOI21X1 AOI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_11661_), .B(_11660_), .C(reset_bF_buf4), .Y(_11521__12_) );
	NAND2X1 NAND2X1_2274 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_13_), .Y(_11662_) );
	NAND2X1 NAND2X1_2275 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf1), .B(_11636__bF_buf1), .Y(_11663_) );
	AOI21X1 AOI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_11663_), .B(_11662_), .C(reset_bF_buf3), .Y(_11521__13_) );
	NAND2X1 NAND2X1_2276 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_14_), .Y(_11664_) );
	NAND2X1 NAND2X1_2277 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf1), .B(_11636__bF_buf0), .Y(_11665_) );
	AOI21X1 AOI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_11665_), .B(_11664_), .C(reset_bF_buf2), .Y(_11521__14_) );
	NAND2X1 NAND2X1_2278 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_15_), .Y(_11666_) );
	NAND2X1 NAND2X1_2279 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf1), .B(_11636__bF_buf4), .Y(_11667_) );
	AOI21X1 AOI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_11667_), .B(_11666_), .C(reset_bF_buf1), .Y(_11521__15_) );
	NAND2X1 NAND2X1_2280 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_16_), .Y(_11668_) );
	NAND2X1 NAND2X1_2281 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_bF_buf1), .B(_11636__bF_buf3), .Y(_11669_) );
	AOI21X1 AOI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_11669_), .B(_11668_), .C(reset_bF_buf0), .Y(_11521__16_) );
	NAND2X1 NAND2X1_2282 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_17_), .Y(_11670_) );
	NAND2X1 NAND2X1_2283 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf1), .B(_11636__bF_buf2), .Y(_11671_) );
	AOI21X1 AOI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_11671_), .B(_11670_), .C(reset_bF_buf10), .Y(_11521__17_) );
	NAND2X1 NAND2X1_2284 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_18_), .Y(_11672_) );
	NAND2X1 NAND2X1_2285 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf0), .B(_11636__bF_buf1), .Y(_11673_) );
	AOI21X1 AOI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_11673_), .B(_11672_), .C(reset_bF_buf9), .Y(_11521__18_) );
	NAND2X1 NAND2X1_2286 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_19_), .Y(_11674_) );
	NAND2X1 NAND2X1_2287 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf3), .B(_11636__bF_buf0), .Y(_11675_) );
	AOI21X1 AOI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_11674_), .C(reset_bF_buf8), .Y(_11521__19_) );
	NAND2X1 NAND2X1_2288 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_20_), .Y(_11676_) );
	NAND2X1 NAND2X1_2289 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf1), .B(_11636__bF_buf4), .Y(_11677_) );
	AOI21X1 AOI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_11677_), .B(_11676_), .C(reset_bF_buf7), .Y(_11521__20_) );
	NAND2X1 NAND2X1_2290 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_21_), .Y(_11678_) );
	NAND2X1 NAND2X1_2291 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf0), .B(_11636__bF_buf3), .Y(_11679_) );
	AOI21X1 AOI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_11679_), .B(_11678_), .C(reset_bF_buf6), .Y(_11521__21_) );
	NAND2X1 NAND2X1_2292 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_22_), .Y(_11680_) );
	NAND2X1 NAND2X1_2293 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf0), .B(_11636__bF_buf2), .Y(_11681_) );
	AOI21X1 AOI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_11681_), .B(_11680_), .C(reset_bF_buf5), .Y(_11521__22_) );
	NAND2X1 NAND2X1_2294 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_23_), .Y(_11682_) );
	NAND2X1 NAND2X1_2295 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_23_), .B(_11636__bF_buf1), .Y(_11683_) );
	AOI21X1 AOI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_11683_), .B(_11682_), .C(reset_bF_buf4), .Y(_11521__23_) );
	NAND2X1 NAND2X1_2296 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_24_), .Y(_11684_) );
	NAND2X1 NAND2X1_2297 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .B(_11636__bF_buf0), .Y(_11685_) );
	AOI21X1 AOI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_11685_), .B(_11684_), .C(reset_bF_buf3), .Y(_11521__24_) );
	NAND2X1 NAND2X1_2298 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_25_), .Y(_11686_) );
	NAND2X1 NAND2X1_2299 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_25_), .B(_11636__bF_buf4), .Y(_11687_) );
	AOI21X1 AOI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_11687_), .B(_11686_), .C(reset_bF_buf2), .Y(_11521__25_) );
	NAND2X1 NAND2X1_2300 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_26_), .Y(_11688_) );
	NAND2X1 NAND2X1_2301 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_26_), .B(_11636__bF_buf3), .Y(_11689_) );
	AOI21X1 AOI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_11689_), .B(_11688_), .C(reset_bF_buf1), .Y(_11521__26_) );
	NAND2X1 NAND2X1_2302 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_27_), .Y(_11690_) );
	NAND2X1 NAND2X1_2303 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_27_), .B(_11636__bF_buf2), .Y(_11691_) );
	AOI21X1 AOI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_11691_), .B(_11690_), .C(reset_bF_buf0), .Y(_11521__27_) );
	NAND2X1 NAND2X1_2304 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_28_), .Y(_11692_) );
	NAND2X1 NAND2X1_2305 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_28_), .B(_11636__bF_buf1), .Y(_11693_) );
	AOI21X1 AOI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_11693_), .B(_11692_), .C(reset_bF_buf10), .Y(_11521__28_) );
	NAND2X1 NAND2X1_2306 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_29_), .Y(_11694_) );
	NAND2X1 NAND2X1_2307 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_29_), .B(_11636__bF_buf0), .Y(_11695_) );
	AOI21X1 AOI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_11695_), .B(_11694_), .C(reset_bF_buf9), .Y(_11521__29_) );
	NAND2X1 NAND2X1_2308 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_30_), .Y(_11696_) );
	NAND2X1 NAND2X1_2309 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_30_), .B(_11636__bF_buf4), .Y(_11697_) );
	AOI21X1 AOI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_11697_), .B(_11696_), .C(reset_bF_buf8), .Y(_11521__30_) );
	NAND2X1 NAND2X1_2310 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(bOperand_frameIn_31_), .Y(_11698_) );
	NAND2X1 NAND2X1_2311 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_B_msb), .B(_11636__bF_buf3), .Y(_11699_) );
	AOI21X1 AOI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_11699_), .B(_11698_), .C(reset_bF_buf7), .Y(_11521__31_) );
	NAND2X1 NAND2X1_2312 ( .gnd(gnd), .vdd(vdd), .A(instructionIn[15]), .B(aLoc_we), .Y(_11700_) );
	INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .Y(_11701_) );
	NAND2X1 NAND2X1_2313 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_0_), .B(_11701_), .Y(_11702_) );
	AOI21X1 AOI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_11702_), .B(_11700_), .C(reset_bF_buf6), .Y(_11518__0_) );
	NAND2X1 NAND2X1_2314 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[16]), .Y(_11703_) );
	NAND2X1 NAND2X1_2315 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .B(_11701_), .Y(_11704_) );
	AOI21X1 AOI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_11704_), .B(_11703_), .C(reset_bF_buf5), .Y(_11518__1_) );
	NAND2X1 NAND2X1_2316 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[17]), .Y(_11705_) );
	NAND2X1 NAND2X1_2317 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_2_), .B(_11701_), .Y(_11706_) );
	AOI21X1 AOI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_11706_), .B(_11705_), .C(reset_bF_buf4), .Y(_11518__2_) );
	NAND2X1 NAND2X1_2318 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[18]), .Y(_11707_) );
	NAND2X1 NAND2X1_2319 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_3_), .B(_11701_), .Y(_11708_) );
	AOI21X1 AOI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_11708_), .B(_11707_), .C(reset_bF_buf3), .Y(_11518__3_) );
	NAND2X1 NAND2X1_2320 ( .gnd(gnd), .vdd(vdd), .A(aLoc_we), .B(instructionIn[19]), .Y(_11709_) );
	NAND2X1 NAND2X1_2321 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(_11701_), .Y(_11710_) );
	AOI21X1 AOI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_11710_), .B(_11709_), .C(reset_bF_buf2), .Y(_11518__4_) );
	NAND2X1 NAND2X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_428__0_), .B(aOperand_we), .Y(_11711_) );
	INVX8 INVX8_47 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .Y(_11712_) );
	NAND2X1 NAND2X1_2323 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf0), .B(_11712__bF_buf4), .Y(_11713_) );
	AOI21X1 AOI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_11713_), .B(_11711_), .C(reset_bF_buf1), .Y(_11519__0_) );
	NAND2X1 NAND2X1_2324 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__1_), .Y(_11714_) );
	NAND2X1 NAND2X1_2325 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf1), .B(_11712__bF_buf3), .Y(_11715_) );
	AOI21X1 AOI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_11715_), .B(_11714_), .C(reset_bF_buf0), .Y(_11519__1_) );
	NAND2X1 NAND2X1_2326 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__2_), .Y(_11716_) );
	NAND2X1 NAND2X1_2327 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf0), .B(_11712__bF_buf2), .Y(_11717_) );
	AOI21X1 AOI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_11717_), .B(_11716_), .C(reset_bF_buf10), .Y(_11519__2_) );
	NAND2X1 NAND2X1_2328 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__3_), .Y(_11718_) );
	NAND2X1 NAND2X1_2329 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(_11712__bF_buf1), .Y(_11719_) );
	AOI21X1 AOI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_11719_), .B(_11718_), .C(reset_bF_buf9), .Y(_11519__3_) );
	NAND2X1 NAND2X1_2330 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__4_), .Y(_11720_) );
	NAND2X1 NAND2X1_2331 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf2), .B(_11712__bF_buf0), .Y(_11721_) );
	AOI21X1 AOI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_11721_), .B(_11720_), .C(reset_bF_buf8), .Y(_11519__4_) );
	NAND2X1 NAND2X1_2332 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__5_), .Y(_11722_) );
	NAND2X1 NAND2X1_2333 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf0), .B(_11712__bF_buf4), .Y(_11723_) );
	AOI21X1 AOI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_11723_), .B(_11722_), .C(reset_bF_buf7), .Y(_11519__5_) );
	NAND2X1 NAND2X1_2334 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__6_), .Y(_11724_) );
	NAND2X1 NAND2X1_2335 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf2), .B(_11712__bF_buf3), .Y(_11725_) );
	AOI21X1 AOI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_11725_), .B(_11724_), .C(reset_bF_buf6), .Y(_11519__6_) );
	NAND2X1 NAND2X1_2336 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__7_), .Y(_11726_) );
	NAND2X1 NAND2X1_2337 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf2), .B(_11712__bF_buf2), .Y(_11727_) );
	AOI21X1 AOI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_11727_), .B(_11726_), .C(reset_bF_buf5), .Y(_11519__7_) );
	NAND2X1 NAND2X1_2338 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__8_), .Y(_11728_) );
	NAND2X1 NAND2X1_2339 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf1), .B(_11712__bF_buf1), .Y(_11729_) );
	AOI21X1 AOI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_11729_), .B(_11728_), .C(reset_bF_buf4), .Y(_11519__8_) );
	NAND2X1 NAND2X1_2340 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__9_), .Y(_11730_) );
	NAND2X1 NAND2X1_2341 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf0), .B(_11712__bF_buf0), .Y(_11731_) );
	AOI21X1 AOI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_11731_), .B(_11730_), .C(reset_bF_buf3), .Y(_11519__9_) );
	NAND2X1 NAND2X1_2342 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__10_), .Y(_11732_) );
	NAND2X1 NAND2X1_2343 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf1), .B(_11712__bF_buf4), .Y(_11733_) );
	AOI21X1 AOI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_11733_), .B(_11732_), .C(reset_bF_buf2), .Y(_11519__10_) );
	NAND2X1 NAND2X1_2344 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__11_), .Y(_11734_) );
	NAND2X1 NAND2X1_2345 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf3), .B(_11712__bF_buf3), .Y(_11735_) );
	AOI21X1 AOI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_11735_), .B(_11734_), .C(reset_bF_buf1), .Y(_11519__11_) );
	NAND2X1 NAND2X1_2346 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__12_), .Y(_11736_) );
	NAND2X1 NAND2X1_2347 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf1), .B(_11712__bF_buf2), .Y(_11737_) );
	AOI21X1 AOI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_11737_), .B(_11736_), .C(reset_bF_buf0), .Y(_11519__12_) );
	NAND2X1 NAND2X1_2348 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__13_), .Y(_11738_) );
	NAND2X1 NAND2X1_2349 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf1), .B(_11712__bF_buf1), .Y(_11739_) );
	AOI21X1 AOI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_11739_), .B(_11738_), .C(reset_bF_buf10), .Y(_11519__13_) );
	NAND2X1 NAND2X1_2350 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__14_), .Y(_11740_) );
	NAND2X1 NAND2X1_2351 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf2), .B(_11712__bF_buf0), .Y(_11741_) );
	AOI21X1 AOI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_11741_), .B(_11740_), .C(reset_bF_buf9), .Y(_11519__14_) );
	NAND2X1 NAND2X1_2352 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__15_), .Y(_11742_) );
	NAND2X1 NAND2X1_2353 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf2), .B(_11712__bF_buf4), .Y(_11743_) );
	AOI21X1 AOI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_11743_), .B(_11742_), .C(reset_bF_buf8), .Y(_11519__15_) );
	NAND2X1 NAND2X1_2354 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__16_), .Y(_11744_) );
	NAND2X1 NAND2X1_2355 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf1), .B(_11712__bF_buf3), .Y(_11745_) );
	AOI21X1 AOI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_11745_), .B(_11744_), .C(reset_bF_buf7), .Y(_11519__16_) );
	NAND2X1 NAND2X1_2356 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__17_), .Y(_11746_) );
	NAND2X1 NAND2X1_2357 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf2), .B(_11712__bF_buf2), .Y(_11747_) );
	AOI21X1 AOI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_11747_), .B(_11746_), .C(reset_bF_buf6), .Y(_11519__17_) );
	NAND2X1 NAND2X1_2358 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__18_), .Y(_11748_) );
	NAND2X1 NAND2X1_2359 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf1), .B(_11712__bF_buf1), .Y(_11749_) );
	AOI21X1 AOI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_11749_), .B(_11748_), .C(reset_bF_buf5), .Y(_11519__18_) );
	NAND2X1 NAND2X1_2360 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__19_), .Y(_11750_) );
	NAND2X1 NAND2X1_2361 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf1), .B(_11712__bF_buf0), .Y(_11751_) );
	AOI21X1 AOI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_11751_), .B(_11750_), .C(reset_bF_buf4), .Y(_11519__19_) );
	NAND2X1 NAND2X1_2362 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__20_), .Y(_11752_) );
	NAND2X1 NAND2X1_2363 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf2), .B(_11712__bF_buf4), .Y(_11753_) );
	AOI21X1 AOI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_11753_), .B(_11752_), .C(reset_bF_buf3), .Y(_11519__20_) );
	NAND2X1 NAND2X1_2364 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__21_), .Y(_11754_) );
	NAND2X1 NAND2X1_2365 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf0), .B(_11712__bF_buf3), .Y(_11755_) );
	AOI21X1 AOI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_11755_), .B(_11754_), .C(reset_bF_buf2), .Y(_11519__21_) );
	NAND2X1 NAND2X1_2366 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__22_), .Y(_11756_) );
	NAND2X1 NAND2X1_2367 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf1), .B(_11712__bF_buf2), .Y(_11757_) );
	AOI21X1 AOI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_11757_), .B(_11756_), .C(reset_bF_buf1), .Y(_11519__22_) );
	NAND2X1 NAND2X1_2368 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__23_), .Y(_11758_) );
	NAND2X1 NAND2X1_2369 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .B(_11712__bF_buf1), .Y(_11759_) );
	AOI21X1 AOI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_11758_), .C(reset_bF_buf0), .Y(_11519__23_) );
	NAND2X1 NAND2X1_2370 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__24_), .Y(_11760_) );
	NAND2X1 NAND2X1_2371 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf3), .B(_11712__bF_buf0), .Y(_11761_) );
	AOI21X1 AOI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_11761_), .B(_11760_), .C(reset_bF_buf10), .Y(_11519__24_) );
	NAND2X1 NAND2X1_2372 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__25_), .Y(_11762_) );
	NAND2X1 NAND2X1_2373 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf0), .B(_11712__bF_buf4), .Y(_11763_) );
	AOI21X1 AOI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_11763_), .B(_11762_), .C(reset_bF_buf9), .Y(_11519__25_) );
	NAND2X1 NAND2X1_2374 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__26_), .Y(_11764_) );
	NAND2X1 NAND2X1_2375 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_26_), .B(_11712__bF_buf3), .Y(_11765_) );
	AOI21X1 AOI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_11765_), .B(_11764_), .C(reset_bF_buf8), .Y(_11519__26_) );
	NAND2X1 NAND2X1_2376 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__27_), .Y(_11766_) );
	NAND2X1 NAND2X1_2377 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_27_), .B(_11712__bF_buf2), .Y(_11767_) );
	AOI21X1 AOI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_11767_), .B(_11766_), .C(reset_bF_buf7), .Y(_11519__27_) );
	NAND2X1 NAND2X1_2378 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__28_), .Y(_11768_) );
	NAND2X1 NAND2X1_2379 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_28_), .B(_11712__bF_buf1), .Y(_11769_) );
	AOI21X1 AOI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_11769_), .B(_11768_), .C(reset_bF_buf6), .Y(_11519__28_) );
	NAND2X1 NAND2X1_2380 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__29_), .Y(_11770_) );
	NAND2X1 NAND2X1_2381 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_29_), .B(_11712__bF_buf0), .Y(_11771_) );
	AOI21X1 AOI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_11771_), .B(_11770_), .C(reset_bF_buf5), .Y(_11519__29_) );
	NAND2X1 NAND2X1_2382 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__30_), .Y(_11772_) );
	NAND2X1 NAND2X1_2383 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .B(_11712__bF_buf4), .Y(_11773_) );
	AOI21X1 AOI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_11773_), .B(_11772_), .C(reset_bF_buf4), .Y(_11519__30_) );
	NAND2X1 NAND2X1_2384 ( .gnd(gnd), .vdd(vdd), .A(aOperand_we), .B(_428__31_), .Y(_11774_) );
	NAND2X1 NAND2X1_2385 ( .gnd(gnd), .vdd(vdd), .A(divider_absoluteValue_A_msb), .B(_11712__bF_buf3), .Y(_11775_) );
	AOI21X1 AOI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_11775_), .B(_11774_), .C(reset_bF_buf3), .Y(_11519__31_) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_11519__0_), .Q(aOperand_frameOut_0_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_11519__1_), .Q(aOperand_frameOut_1_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_11519__2_), .Q(aOperand_frameOut_2_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_11519__3_), .Q(aOperand_frameOut_3_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_11519__4_), .Q(aOperand_frameOut_4_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_11519__5_), .Q(aOperand_frameOut_5_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_11519__6_), .Q(aOperand_frameOut_6_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_11519__7_), .Q(aOperand_frameOut_7_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_11519__8_), .Q(aOperand_frameOut_8_) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_11519__9_), .Q(aOperand_frameOut_9_) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_11519__10_), .Q(aOperand_frameOut_10_) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_11519__11_), .Q(aOperand_frameOut_11_) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_11519__12_), .Q(aOperand_frameOut_12_) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_11519__13_), .Q(aOperand_frameOut_13_) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_11519__14_), .Q(aOperand_frameOut_14_) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_11519__15_), .Q(aOperand_frameOut_15_) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_11519__16_), .Q(aOperand_frameOut_16_) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_11519__17_), .Q(aOperand_frameOut_17_) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_11519__18_), .Q(aOperand_frameOut_18_) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_11519__19_), .Q(aOperand_frameOut_19_) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_11519__20_), .Q(aOperand_frameOut_20_) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_11519__21_), .Q(aOperand_frameOut_21_) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_11519__22_), .Q(aOperand_frameOut_22_) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_11519__23_), .Q(aOperand_frameOut_23_) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_11519__24_), .Q(aOperand_frameOut_24_) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_11519__25_), .Q(aOperand_frameOut_25_) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_11519__26_), .Q(aOperand_frameOut_26_) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_11519__27_), .Q(aOperand_frameOut_27_) );
	DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_11519__28_), .Q(aOperand_frameOut_28_) );
	DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_11519__29_), .Q(aOperand_frameOut_29_) );
	DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_11519__30_), .Q(aOperand_frameOut_30_) );
	DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_11519__31_), .Q(divider_absoluteValue_A_msb) );
	DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_11518__0_), .Q(aLoc_frameOut_0_) );
	DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_11518__1_), .Q(aLoc_frameOut_1_) );
	DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_11518__2_), .Q(aLoc_frameOut_2_) );
	DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_11518__3_), .Q(aLoc_frameOut_3_) );
	DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_11518__4_), .Q(aLoc_frameOut_4_) );
	DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_11521__0_), .Q(adder_bOperand_0_) );
	DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_11521__1_), .Q(adder_bOperand_1_) );
	DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_11521__2_), .Q(adder_bOperand_2_) );
	DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_11521__3_), .Q(adder_bOperand_3_) );
	DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_11521__4_), .Q(adder_bOperand_4_) );
	DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_11521__5_), .Q(adder_bOperand_5_) );
	DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_11521__6_), .Q(adder_bOperand_6_) );
	DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_11521__7_), .Q(adder_bOperand_7_) );
	DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_11521__8_), .Q(adder_bOperand_8_) );
	DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_11521__9_), .Q(adder_bOperand_9_) );
	DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_11521__10_), .Q(adder_bOperand_10_) );
	DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_11521__11_), .Q(adder_bOperand_11_) );
	DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_11521__12_), .Q(adder_bOperand_12_) );
	DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_11521__13_), .Q(adder_bOperand_13_) );
	DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_11521__14_), .Q(adder_bOperand_14_) );
	DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_11521__15_), .Q(adder_bOperand_15_) );
	DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_11521__16_), .Q(adder_bOperand_16_) );
	DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_11521__17_), .Q(adder_bOperand_17_) );
	DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_11521__18_), .Q(adder_bOperand_18_) );
	DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_11521__19_), .Q(adder_bOperand_19_) );
	DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_11521__20_), .Q(adder_bOperand_20_) );
	DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_11521__21_), .Q(adder_bOperand_21_) );
	DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_11521__22_), .Q(adder_bOperand_22_) );
	DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_11521__23_), .Q(adder_bOperand_23_) );
	DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_11521__24_), .Q(adder_bOperand_24_) );
	DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_11521__25_), .Q(adder_bOperand_25_) );
	DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_11521__26_), .Q(adder_bOperand_26_) );
	DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_11521__27_), .Q(adder_bOperand_27_) );
	DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_11521__28_), .Q(adder_bOperand_28_) );
	DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_11521__29_), .Q(adder_bOperand_29_) );
	DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_11521__30_), .Q(adder_bOperand_30_) );
	DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_11521__31_), .Q(divider_absoluteValue_B_msb) );
	DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_11520__0_), .Q(bLoc_frameOut_0_) );
	DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_11520__1_), .Q(bLoc_frameOut_1_) );
	DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_11520__2_), .Q(bLoc_frameOut_2_) );
	DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_11520__3_), .Q(bLoc_frameOut_3_) );
	DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_11520__4_), .Q(bLoc_frameOut_4_) );
	DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_11523__0_), .Q(immediateVal_frameOut_0_) );
	DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_11523__1_), .Q(immediateVal_frameOut_1_) );
	DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_11523__2_), .Q(immediateVal_frameOut_2_) );
	DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_11523__3_), .Q(immediateVal_frameOut_3_) );
	DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_11523__4_), .Q(immediateVal_frameOut_4_) );
	DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_11523__5_), .Q(immediateVal_frameOut_5_) );
	DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_11523__6_), .Q(immediateVal_frameOut_6_) );
	DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_11523__7_), .Q(immediateVal_frameOut_7_) );
	DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_11523__8_), .Q(immediateVal_frameOut_8_) );
	DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_11523__9_), .Q(immediateVal_frameOut_9_) );
	DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_11523__10_), .Q(immediateVal_frameOut_10_) );
	DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_11523__11_), .Q(immediateVal_frameOut_11_) );
	DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_11523__12_), .Q(immediateVal_frameOut_12_) );
	DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_11523__13_), .Q(immediateVal_frameOut_13_) );
	DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_11523__14_), .Q(immediateVal_frameOut_14_) );
	DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_11523__15_), .Q(immediateVal_frameOut_15_) );
	DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_11523__16_), .Q(immediateVal_frameOut_16_) );
	DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_11523__17_), .Q(immediateVal_frameOut_17_) );
	DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_11523__18_), .Q(immediateVal_frameOut_18_) );
	DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_11523__19_), .Q(immediateVal_frameOut_19_) );
	DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_11523__20_), .Q(immediateVal_frameOut_20_) );
	DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_11523__21_), .Q(immediateVal_frameOut_21_) );
	DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_11523__22_), .Q(immediateVal_frameOut_22_) );
	DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_11523__23_), .Q(immediateVal_frameOut_23_) );
	DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_11523__24_), .Q(immediateVal_frameOut_24_) );
	DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_11523__25_), .Q(immediateVal_frameOut_25_) );
	DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_11523__26_), .Q(immediateVal_frameOut_26_) );
	DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_11523__27_), .Q(immediateVal_frameOut_27_) );
	DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_11523__28_), .Q(immediateVal_frameOut_28_) );
	DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_11523__29_), .Q(immediateVal_frameOut_29_) );
	DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_11523__30_), .Q(immediateVal_frameOut_30_) );
	DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_11523__31_), .Q(immediateVal_frameOut_31_) );
	DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_11522_), .Q(immediateSelect_frameOut) );
	DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_11526_), .Q(comparator_unsignedEn) );
	DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_11525_), .Q(adder_subtract) );
	DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_11524__0_), .Q(instructionFrame_resultSelect_out_0_) );
	DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_11524__1_), .Q(instructionFrame_resultSelect_out_1_) );
	DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_11524__2_), .Q(instructionFrame_resultSelect_out_2_) );
	DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_11528__0_), .Q(instructionFrame_writeSelect_out_0_) );
	DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_11528__1_), .Q(instructionFrame_writeSelect_out_1_) );
	DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_11528__2_), .Q(instructionFrame_writeSelect_out_2_) );
	DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_11528__3_), .Q(instructionFrame_writeSelect_out_3_) );
	DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_11528__4_), .Q(instructionFrame_writeSelect_out_4_) );
	DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_11527_), .Q(instructionFrame_writeEnable_out) );
	INVX8 INVX8_48 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .Y(_17295_) );
	INVX8 INVX8_49 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf4), .Y(_17306_) );
	NOR2X1 NOR2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf4), .B(_17306__bF_buf3), .Y(mulOut_0_) );
	INVX8 INVX8_50 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf4), .Y(_11776_) );
	NOR2X1 NOR2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf2), .B(_11776__bF_buf3), .Y(_11797_) );
	NAND2X1 NAND2X1_2386 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_1_bF_buf0), .Y(_11798_) );
	INVX1 INVX1_1639 ( .gnd(gnd), .vdd(vdd), .A(_11798_), .Y(_11809_) );
	AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_11797_), .B(_11809_), .Y(_11820_) );
	NOR2X1 NOR2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_11809_), .B(_11797_), .Y(_11831_) );
	NOR2X1 NOR2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_11831_), .B(_11820_), .Y(mulOut_1_) );
	NAND2X1 NAND2X1_2387 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf3), .B(adder_bOperand_2_bF_buf0), .Y(_11852_) );
	NAND2X1 NAND2X1_2388 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf3), .B(aOperand_frameOut_2_bF_buf4), .Y(_11863_) );
	INVX8 INVX8_51 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf5), .Y(_11874_) );
	NAND2X1 NAND2X1_2389 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_2_bF_buf3), .Y(_11885_) );
	OAI21X1 OAI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_11776__bF_buf2), .C(_11885_), .Y(_11906_) );
	OAI21X1 OAI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_11798_), .B(_11863_), .C(_11906_), .Y(_11917_) );
	XOR2X1 XOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_11917_), .B(_11852_), .Y(_11918_) );
	NAND2X1 NAND2X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_11820_), .B(_11918_), .Y(_11929_) );
	INVX1 INVX1_1640 ( .gnd(gnd), .vdd(vdd), .A(_11929_), .Y(_11939_) );
	NOR2X1 NOR2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_11820_), .B(_11918_), .Y(_11950_) );
	NOR2X1 NOR2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_11950_), .B(_11939_), .Y(mulOut_2_) );
	INVX8 INVX8_52 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf2), .Y(_11971_) );
	NOR2X1 NOR2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf1), .B(_11971__bF_buf3), .Y(_11982_) );
	INVX1 INVX1_1641 ( .gnd(gnd), .vdd(vdd), .A(_11863_), .Y(_11993_) );
	NOR2X1 NOR2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_11852_), .B(_11917_), .Y(_12004_) );
	AOI21X1 AOI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_11809_), .B(_11993_), .C(_12004_), .Y(_12015_) );
	NAND2X1 NAND2X1_2391 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf4), .B(adder_bOperand_2_bF_buf5), .Y(_12026_) );
	NAND2X1 NAND2X1_2392 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .B(aOperand_frameOut_3_bF_buf0), .Y(_12037_) );
	INVX8 INVX8_53 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf4), .Y(_12048_) );
	OAI21X1 OAI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf3), .B(_12048_), .C(_11863_), .Y(_12059_) );
	OAI21X1 OAI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_11885_), .B(_12037_), .C(_12059_), .Y(_12070_) );
	OR2X2 OR2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_12070_), .B(_12026_), .Y(_12081_) );
	INVX8 INVX8_54 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .Y(_12092_) );
	OAI21X1 OAI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_12092_), .C(_12070_), .Y(_12103_) );
	NAND2X1 NAND2X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_12103_), .B(_12081_), .Y(_12114_) );
	NOR2X1 NOR2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_12015_), .B(_12114_), .Y(_12124_) );
	AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_12114_), .B(_12015_), .Y(_12135_) );
	NOR2X1 NOR2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_12124_), .B(_12135_), .Y(_12146_) );
	NAND2X1 NAND2X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_11982_), .B(_12146_), .Y(_12157_) );
	INVX1 INVX1_1642 ( .gnd(gnd), .vdd(vdd), .A(_11982_), .Y(_12178_) );
	OAI21X1 OAI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_12124_), .B(_12135_), .C(_12178_), .Y(_12179_) );
	AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_12157_), .B(_12179_), .Y(_12190_) );
	NAND2X1 NAND2X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_11939_), .B(_12190_), .Y(_12201_) );
	INVX1 INVX1_1643 ( .gnd(gnd), .vdd(vdd), .A(_12201_), .Y(_12212_) );
	NOR2X1 NOR2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_11939_), .B(_12190_), .Y(_12223_) );
	NOR2X1 NOR2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_12223_), .B(_12212_), .Y(mulOut_3_) );
	OAI21X1 OAI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_12015_), .B(_12114_), .C(_12157_), .Y(_12244_) );
	NAND2X1 NAND2X1_2396 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf3), .B(adder_bOperand_4_bF_buf3), .Y(_12255_) );
	INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf2), .Y(_12266_) );
	OAI22X1 OAI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf0), .B(_12266_), .C(_11874_), .D(_11971__bF_buf2), .Y(_12277_) );
	OAI21X1 OAI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_12255_), .B(_12178_), .C(_12277_), .Y(_12288_) );
	OAI21X1 OAI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_11885_), .B(_12037_), .C(_12081_), .Y(_12299_) );
	INVX8 INVX8_55 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf2), .Y(_12310_) );
	NOR2X1 NOR2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf3), .B(_12092_), .Y(_12320_) );
	NAND2X1 NAND2X1_2397 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_3_bF_buf3), .Y(_12341_) );
	NAND2X1 NAND2X1_2398 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf1), .B(aOperand_frameOut_4_bF_buf1), .Y(_12352_) );
	INVX8 INVX8_56 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf0), .Y(_12353_) );
	OAI21X1 OAI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf2), .B(_12353__bF_buf3), .C(_12037_), .Y(_12364_) );
	OAI21X1 OAI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_12341_), .B(_12352_), .C(_12364_), .Y(_12375_) );
	XNOR2X1 XNOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12320_), .Y(_12386_) );
	NAND2X1 NAND2X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_12386_), .B(_12299_), .Y(_12397_) );
	INVX1 INVX1_1644 ( .gnd(gnd), .vdd(vdd), .A(_12341_), .Y(_12408_) );
	NOR2X1 NOR2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_12026_), .B(_12070_), .Y(_12419_) );
	AOI21X1 AOI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_11993_), .B(_12408_), .C(_12419_), .Y(_12430_) );
	XOR2X1 XOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12320_), .Y(_12441_) );
	NAND2X1 NAND2X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_12441_), .B(_12430_), .Y(_12452_) );
	NAND2X1 NAND2X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_12452_), .B(_12397_), .Y(_12463_) );
	NOR2X1 NOR2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_12288_), .B(_12463_), .Y(_12474_) );
	INVX1 INVX1_1645 ( .gnd(gnd), .vdd(vdd), .A(_12288_), .Y(_12485_) );
	AOI21X1 AOI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_12397_), .B(_12452_), .C(_12485_), .Y(_12496_) );
	OAI21X1 OAI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_12474_), .B(_12496_), .C(_12244_), .Y(_12507_) );
	INVX1 INVX1_1646 ( .gnd(gnd), .vdd(vdd), .A(_12244_), .Y(_12518_) );
	NOR2X1 NOR2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_12496_), .B(_12474_), .Y(_12529_) );
	NAND2X1 NAND2X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .B(_12518_), .Y(_12540_) );
	AOI21X1 AOI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_12540_), .B(_12507_), .C(_12201_), .Y(_12551_) );
	NAND2X1 NAND2X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_12507_), .B(_12540_), .Y(_12561_) );
	NOR2X1 NOR2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_12212_), .B(_12561_), .Y(_12572_) );
	NOR2X1 NOR2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_12551_), .B(_12572_), .Y(mulOut_4_) );
	NAND2X1 NAND2X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .B(_12244_), .Y(_12593_) );
	INVX1 INVX1_1647 ( .gnd(gnd), .vdd(vdd), .A(_12593_), .Y(_12614_) );
	OR2X2 OR2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_12178_), .B(_12255_), .Y(_12615_) );
	INVX1 INVX1_1648 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .Y(_12626_) );
	NOR2X1 NOR2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_12441_), .B(_12430_), .Y(_12637_) );
	AOI21X1 AOI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_12485_), .B(_12452_), .C(_12637_), .Y(_12648_) );
	NAND2X1 NAND2X1_2405 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf2), .B(adder_bOperand_5_bF_buf0), .Y(_12659_) );
	NAND2X1 NAND2X1_2406 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf1), .B(adder_bOperand_3_bF_buf1), .Y(_12670_) );
	XOR2X1 XOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_12255_), .B(_12670_), .Y(_12681_) );
	XNOR2X1 XNOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_12681_), .B(_12659_), .Y(_12692_) );
	INVX1 INVX1_1649 ( .gnd(gnd), .vdd(vdd), .A(_12352_), .Y(_12703_) );
	AOI22X1 AOI22X1_269 ( .gnd(gnd), .vdd(vdd), .A(_12408_), .B(_12703_), .C(_12320_), .D(_12364_), .Y(_12714_) );
	INVX1 INVX1_1650 ( .gnd(gnd), .vdd(vdd), .A(_12714_), .Y(_12725_) );
	NOR2X1 NOR2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12048_), .Y(_12736_) );
	NAND2X1 NAND2X1_2407 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(aOperand_frameOut_5_bF_buf4), .Y(_12747_) );
	NOR2X1 NOR2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_12352_), .B(_12747_), .Y(_12758_) );
	INVX1 INVX1_1651 ( .gnd(gnd), .vdd(vdd), .A(_12758_), .Y(_12769_) );
	INVX8 INVX8_57 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf3), .Y(_12780_) );
	OAI21X1 OAI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf1), .B(_12780_), .C(_12352_), .Y(_12790_) );
	NAND3X1 NAND3X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_12736_), .B(_12790_), .C(_12769_), .Y(_12801_) );
	NAND2X1 NAND2X1_2408 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .B(aOperand_frameOut_4_bF_buf4), .Y(_12812_) );
	NAND2X1 NAND2X1_2409 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf0), .B(aOperand_frameOut_5_bF_buf2), .Y(_12833_) );
	OAI21X1 OAI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_12812_), .B(_12833_), .C(_12790_), .Y(_12844_) );
	OAI21X1 OAI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12048_), .C(_12844_), .Y(_12845_) );
	NAND3X1 NAND3X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_12801_), .B(_12845_), .C(_12725_), .Y(_12866_) );
	NAND2X1 NAND2X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_12801_), .B(_12845_), .Y(_12867_) );
	NAND2X1 NAND2X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_12714_), .B(_12867_), .Y(_12878_) );
	NAND3X1 NAND3X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_12692_), .B(_12866_), .C(_12878_), .Y(_12889_) );
	INVX1 INVX1_1652 ( .gnd(gnd), .vdd(vdd), .A(_12889_), .Y(_12900_) );
	AOI21X1 AOI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_12878_), .B(_12866_), .C(_12692_), .Y(_12911_) );
	NOR3X1 NOR3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_12911_), .B(_12648_), .C(_12900_), .Y(_12922_) );
	INVX1 INVX1_1653 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .Y(_12933_) );
	OAI21X1 OAI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_12911_), .B(_12900_), .C(_12648_), .Y(_12944_) );
	NAND3X1 NAND3X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_12626_), .B(_12944_), .C(_12933_), .Y(_12955_) );
	INVX1 INVX1_1654 ( .gnd(gnd), .vdd(vdd), .A(_12944_), .Y(_12966_) );
	OAI21X1 OAI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .B(_12966_), .C(_12615_), .Y(_12977_) );
	NAND3X1 NAND3X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_12955_), .B(_12977_), .C(_12614_), .Y(_12988_) );
	NAND3X1 NAND3X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .B(_12944_), .C(_12933_), .Y(_12999_) );
	OAI21X1 OAI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_12922_), .B(_12966_), .C(_12626_), .Y(_13010_) );
	NAND3X1 NAND3X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_12593_), .B(_13010_), .C(_12999_), .Y(_13021_) );
	NAND3X1 NAND3X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_12988_), .B(_13021_), .C(_12551_), .Y(_13032_) );
	INVX1 INVX1_1655 ( .gnd(gnd), .vdd(vdd), .A(_13032_), .Y(_13043_) );
	AOI21X1 AOI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_12988_), .B(_13021_), .C(_12551_), .Y(_13054_) );
	NOR2X1 NOR2X1_784 ( .gnd(gnd), .vdd(vdd), .A(_13054_), .B(_13043_), .Y(mulOut_5_) );
	OAI21X1 OAI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .B(_12966_), .C(_12933_), .Y(_13074_) );
	NAND2X1 NAND2X1_2412 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf1), .B(adder_bOperand_6_bF_buf2), .Y(_13085_) );
	INVX1 INVX1_1656 ( .gnd(gnd), .vdd(vdd), .A(_13085_), .Y(_13096_) );
	NAND3X1 NAND3X1_2331 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf0), .B(adder_bOperand_5_bF_buf4), .C(_12681_), .Y(_13107_) );
	OAI21X1 OAI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_12255_), .B(_12670_), .C(_13107_), .Y(_13118_) );
	XNOR2X1 XNOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_13118_), .B(_13096_), .Y(_13129_) );
	XOR2X1 XOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_12681_), .B(_12659_), .Y(_13140_) );
	AOI21X1 AOI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_12845_), .B(_12801_), .C(_12725_), .Y(_13151_) );
	OAI21X1 OAI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13140_), .C(_12866_), .Y(_13162_) );
	NAND2X1 NAND2X1_2413 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf2), .B(adder_bOperand_5_bF_buf3), .Y(_13173_) );
	NAND2X1 NAND2X1_2414 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .B(adder_bOperand_4_bF_buf1), .Y(_13184_) );
	NAND2X1 NAND2X1_2415 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(adder_bOperand_3_bF_buf0), .Y(_13195_) );
	OAI21X1 OAI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf2), .B(_12266_), .C(_13195_), .Y(_13206_) );
	OAI21X1 OAI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_12670_), .B(_13184_), .C(_13206_), .Y(_13217_) );
	XOR2X1 XOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .B(_13173_), .Y(_13228_) );
	AOI21X1 AOI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_12790_), .B(_12736_), .C(_12758_), .Y(_13239_) );
	INVX1 INVX1_1657 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .Y(_13250_) );
	NOR2X1 NOR2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12353__bF_buf2), .Y(_13261_) );
	INVX1 INVX1_1658 ( .gnd(gnd), .vdd(vdd), .A(_13261_), .Y(_13272_) );
	NAND2X1 NAND2X1_2416 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf6), .B(aOperand_frameOut_6_bF_buf1), .Y(_13283_) );
	INVX8 INVX8_58 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf0), .Y(_13294_) );
	OAI21X1 OAI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf0), .B(_13294__bF_buf3), .C(_12833_), .Y(_13305_) );
	OAI21X1 OAI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_12747_), .B(_13283_), .C(_13305_), .Y(_13316_) );
	OR2X2 OR2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_13316_), .B(_13272_), .Y(_13326_) );
	OAI21X1 OAI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12353__bF_buf1), .C(_13316_), .Y(_13337_) );
	NAND3X1 NAND3X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_13337_), .B(_13250_), .C(_13326_), .Y(_13348_) );
	NOR2X1 NOR2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_13272_), .B(_13316_), .Y(_13359_) );
	INVX1 INVX1_1659 ( .gnd(gnd), .vdd(vdd), .A(_12747_), .Y(_13370_) );
	INVX1 INVX1_1660 ( .gnd(gnd), .vdd(vdd), .A(_13283_), .Y(_13381_) );
	NAND2X1 NAND2X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_13370_), .B(_13381_), .Y(_13392_) );
	AOI21X1 AOI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_13392_), .B(_13305_), .C(_13261_), .Y(_13403_) );
	OAI21X1 OAI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13359_), .C(_13239_), .Y(_13414_) );
	NAND3X1 NAND3X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_13228_), .B(_13414_), .C(_13348_), .Y(_13425_) );
	INVX8 INVX8_59 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf2), .Y(_13436_) );
	OAI21X1 OAI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_13436__bF_buf3), .C(_13217_), .Y(_13447_) );
	OR2X2 OR2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_13217_), .B(_13173_), .Y(_13458_) );
	NAND2X1 NAND2X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_13447_), .B(_13458_), .Y(_13469_) );
	OAI21X1 OAI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_13403_), .B(_13359_), .C(_13250_), .Y(_13480_) );
	NAND3X1 NAND3X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .B(_13337_), .C(_13326_), .Y(_13491_) );
	NAND3X1 NAND3X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_13469_), .B(_13480_), .C(_13491_), .Y(_13502_) );
	NAND3X1 NAND3X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_13425_), .B(_13502_), .C(_13162_), .Y(_13513_) );
	INVX1 INVX1_1661 ( .gnd(gnd), .vdd(vdd), .A(_13162_), .Y(_13524_) );
	NAND2X1 NAND2X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_13425_), .B(_13502_), .Y(_13535_) );
	NAND2X1 NAND2X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_13524_), .B(_13535_), .Y(_13546_) );
	NAND2X1 NAND2X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_13513_), .B(_13546_), .Y(_13557_) );
	NOR2X1 NOR2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_13129_), .B(_13557_), .Y(_13568_) );
	INVX1 INVX1_1662 ( .gnd(gnd), .vdd(vdd), .A(_13129_), .Y(_13579_) );
	AOI21X1 AOI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_13546_), .B(_13513_), .C(_13579_), .Y(_13600_) );
	OAI21X1 OAI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_13568_), .B(_13600_), .C(_13074_), .Y(_13601_) );
	AOI21X1 AOI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_12626_), .B(_12944_), .C(_12922_), .Y(_13621_) );
	OR2X2 OR2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_13557_), .B(_13129_), .Y(_13622_) );
	INVX1 INVX1_1663 ( .gnd(gnd), .vdd(vdd), .A(_13600_), .Y(_13633_) );
	NAND3X1 NAND3X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_13621_), .B(_13633_), .C(_13622_), .Y(_13644_) );
	NAND2X1 NAND2X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_13644_), .B(_13601_), .Y(_13655_) );
	NAND2X1 NAND2X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_12988_), .B(_13655_), .Y(_13666_) );
	AOI21X1 AOI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_12999_), .B(_13010_), .C(_12593_), .Y(_13677_) );
	NAND3X1 NAND3X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_13601_), .B(_13644_), .C(_13677_), .Y(_13688_) );
	AOI21X1 AOI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_13666_), .B(_13688_), .C(_13032_), .Y(_13699_) );
	NAND2X1 NAND2X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_13688_), .B(_13666_), .Y(_13710_) );
	NOR2X1 NOR2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_13043_), .B(_13710_), .Y(_13721_) );
	NOR2X1 NOR2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_13699_), .B(_13721_), .Y(mulOut_6_) );
	NAND3X1 NAND3X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_13633_), .B(_13622_), .C(_13074_), .Y(_13742_) );
	NAND2X1 NAND2X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_13096_), .B(_13118_), .Y(_13753_) );
	INVX1 INVX1_1664 ( .gnd(gnd), .vdd(vdd), .A(_13753_), .Y(_13764_) );
	AOI21X1 AOI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_13502_), .B(_13425_), .C(_13162_), .Y(_13775_) );
	OAI21X1 OAI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_13129_), .B(_13775_), .C(_13513_), .Y(_13786_) );
	NAND2X1 NAND2X1_2426 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf1), .B(adder_bOperand_7_bF_buf3), .Y(_13797_) );
	NOR2X1 NOR2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_13085_), .B(_13797_), .Y(_13808_) );
	INVX1 INVX1_1665 ( .gnd(gnd), .vdd(vdd), .A(_13808_), .Y(_13819_) );
	INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf2), .Y(_13830_) );
	NAND2X1 NAND2X1_2427 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf0), .B(adder_bOperand_6_bF_buf1), .Y(_13841_) );
	OAI21X1 OAI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf3), .B(_13830_), .C(_13841_), .Y(_13852_) );
	AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_13819_), .B(_13852_), .Y(_13863_) );
	OAI21X1 OAI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_12670_), .B(_13184_), .C(_13458_), .Y(_13874_) );
	XNOR2X1 XNOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_13874_), .B(_13863_), .Y(_13885_) );
	INVX1 INVX1_1666 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .Y(_13896_) );
	AOI21X1 AOI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_13326_), .B(_13337_), .C(_13250_), .Y(_13906_) );
	OAI21X1 OAI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_13469_), .B(_13906_), .C(_13348_), .Y(_13917_) );
	NOR2X1 NOR2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf1), .B(_13436__bF_buf2), .Y(_13928_) );
	NAND2X1 NAND2X1_2428 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .B(adder_bOperand_4_bF_buf0), .Y(_13939_) );
	OAI21X1 OAI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf1), .B(_12353__bF_buf0), .C(_13184_), .Y(_13950_) );
	OAI21X1 OAI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_13195_), .B(_13939_), .C(_13950_), .Y(_13961_) );
	XNOR2X1 XNOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_13961_), .B(_13928_), .Y(_13972_) );
	AOI22X1 AOI22X1_270 ( .gnd(gnd), .vdd(vdd), .A(_13370_), .B(_13381_), .C(_13261_), .D(_13305_), .Y(_13983_) );
	INVX1 INVX1_1667 ( .gnd(gnd), .vdd(vdd), .A(_13983_), .Y(_13994_) );
	NOR2X1 NOR2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12780_), .Y(_14005_) );
	NAND2X1 NAND2X1_2429 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(aOperand_frameOut_7_bF_buf1), .Y(_14016_) );
	NOR2X1 NOR2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_13283_), .B(_14016_), .Y(_14037_) );
	INVX1 INVX1_1668 ( .gnd(gnd), .vdd(vdd), .A(_14037_), .Y(_14048_) );
	INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf0), .Y(_14049_) );
	OAI21X1 OAI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf4), .B(_14049_), .C(_13283_), .Y(_14060_) );
	NAND3X1 NAND3X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_14005_), .B(_14060_), .C(_14048_), .Y(_14071_) );
	NAND2X1 NAND2X1_2430 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .B(aOperand_frameOut_6_bF_buf4), .Y(_14082_) );
	NAND2X1 NAND2X1_2431 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(aOperand_frameOut_7_bF_buf4), .Y(_14093_) );
	OAI21X1 OAI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_14082_), .B(_14093_), .C(_14060_), .Y(_14104_) );
	OAI21X1 OAI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_12780_), .C(_14104_), .Y(_14115_) );
	NAND3X1 NAND3X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_14071_), .B(_14115_), .C(_13994_), .Y(_14126_) );
	INVX1 INVX1_1669 ( .gnd(gnd), .vdd(vdd), .A(_14005_), .Y(_14137_) );
	NOR2X1 NOR2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_14137_), .B(_14104_), .Y(_14148_) );
	AOI21X1 AOI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_14048_), .B(_14060_), .C(_14005_), .Y(_14159_) );
	OAI21X1 OAI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_14148_), .B(_14159_), .C(_13983_), .Y(_14170_) );
	NAND3X1 NAND3X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_14126_), .B(_13972_), .C(_14170_), .Y(_14181_) );
	XOR2X1 XOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_13961_), .B(_13928_), .Y(_14192_) );
	OAI21X1 OAI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_14148_), .B(_14159_), .C(_13994_), .Y(_14203_) );
	NAND3X1 NAND3X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_13983_), .B(_14071_), .C(_14115_), .Y(_14214_) );
	NAND3X1 NAND3X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_14192_), .B(_14214_), .C(_14203_), .Y(_14225_) );
	NAND3X1 NAND3X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_14181_), .B(_14225_), .C(_13917_), .Y(_14235_) );
	NOR3X1 NOR3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_13239_), .B(_13403_), .C(_13359_), .Y(_14246_) );
	AOI21X1 AOI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_13228_), .B(_13414_), .C(_14246_), .Y(_14257_) );
	AOI21X1 AOI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_14203_), .B(_14214_), .C(_14192_), .Y(_14268_) );
	AOI21X1 AOI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_14170_), .B(_14126_), .C(_13972_), .Y(_14279_) );
	OAI21X1 OAI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(_14279_), .C(_14257_), .Y(_14290_) );
	NAND3X1 NAND3X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_14235_), .B(_14290_), .C(_13896_), .Y(_14301_) );
	OAI21X1 OAI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(_14279_), .C(_13917_), .Y(_14312_) );
	NAND3X1 NAND3X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_14181_), .B(_14225_), .C(_14257_), .Y(_14323_) );
	NAND3X1 NAND3X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .B(_14323_), .C(_14312_), .Y(_14334_) );
	NAND3X1 NAND3X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_13786_), .B(_14334_), .C(_14301_), .Y(_14345_) );
	INVX1 INVX1_1670 ( .gnd(gnd), .vdd(vdd), .A(_13786_), .Y(_14356_) );
	AOI21X1 AOI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_14312_), .B(_14323_), .C(_13885_), .Y(_14367_) );
	AOI21X1 AOI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_14290_), .B(_14235_), .C(_13896_), .Y(_14378_) );
	OAI21X1 OAI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_14367_), .B(_14378_), .C(_14356_), .Y(_14389_) );
	NAND3X1 NAND3X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_14345_), .C(_14389_), .Y(_14400_) );
	OAI21X1 OAI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_14367_), .B(_14378_), .C(_13786_), .Y(_14411_) );
	NAND3X1 NAND3X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_14301_), .B(_14334_), .C(_14356_), .Y(_14422_) );
	NAND3X1 NAND3X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_13753_), .B(_14411_), .C(_14422_), .Y(_14433_) );
	NAND3X1 NAND3X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_13742_), .B(_14400_), .C(_14433_), .Y(_14444_) );
	NOR3X1 NOR3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_13600_), .B(_13621_), .C(_13568_), .Y(_14455_) );
	NAND3X1 NAND3X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_13753_), .B(_14345_), .C(_14389_), .Y(_14466_) );
	NAND3X1 NAND3X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_14411_), .C(_14422_), .Y(_14477_) );
	NAND3X1 NAND3X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_14455_), .B(_14466_), .C(_14477_), .Y(_14498_) );
	NAND2X1 NAND2X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_14444_), .B(_14498_), .Y(_14499_) );
	AOI21X1 AOI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_13601_), .B(_13644_), .C(_12988_), .Y(_14510_) );
	NOR2X1 NOR2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_14510_), .B(_13699_), .Y(_14521_) );
	XNOR2X1 XNOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_14521_), .B(_14499_), .Y(mulOut_7_) );
	NAND2X1 NAND2X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_14499_), .B(_13699_), .Y(_14541_) );
	NAND3X1 NAND3X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_14455_), .B(_14400_), .C(_14433_), .Y(_14552_) );
	NAND3X1 NAND3X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_13742_), .B(_14466_), .C(_14477_), .Y(_14563_) );
	NAND3X1 NAND3X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_14552_), .B(_14563_), .C(_14510_), .Y(_14574_) );
	AOI21X1 AOI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_14477_), .B(_14466_), .C(_13742_), .Y(_14585_) );
	AOI21X1 AOI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_14301_), .B(_14334_), .C(_13786_), .Y(_14596_) );
	OAI21X1 OAI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_13753_), .B(_14596_), .C(_14345_), .Y(_14607_) );
	NAND2X1 NAND2X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_13863_), .B(_13874_), .Y(_14618_) );
	INVX1 INVX1_1671 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .Y(_14629_) );
	AOI21X1 AOI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_14181_), .B(_14225_), .C(_13917_), .Y(_14640_) );
	OAI21X1 OAI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_13885_), .B(_14640_), .C(_14235_), .Y(_14651_) );
	NAND2X1 NAND2X1_2435 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf4), .B(adder_bOperand_8_bF_buf0), .Y(_14662_) );
	NAND2X1 NAND2X1_2436 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf0), .B(adder_bOperand_7_bF_buf1), .Y(_14673_) );
	INVX8 INVX8_60 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf0), .Y(_14684_) );
	OAI21X1 OAI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf0), .B(_14684__bF_buf3), .C(_13797_), .Y(_14695_) );
	OAI21X1 OAI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_13841_), .B(_14673_), .C(_14695_), .Y(_14706_) );
	OR2X2 OR2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_14706_), .B(_14662_), .Y(_14717_) );
	INVX8 INVX8_61 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf4), .Y(_14728_) );
	OAI21X1 OAI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf2), .B(_14728__bF_buf3), .C(_14706_), .Y(_14749_) );
	NAND2X1 NAND2X1_2437 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf5), .B(aOperand_frameOut_4_bF_buf2), .Y(_14760_) );
	NOR2X1 NOR2X1_796 ( .gnd(gnd), .vdd(vdd), .A(_13184_), .B(_14760_), .Y(_14761_) );
	AOI21X1 AOI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_13950_), .B(_13928_), .C(_14761_), .Y(_14772_) );
	INVX1 INVX1_1672 ( .gnd(gnd), .vdd(vdd), .A(_14772_), .Y(_14783_) );
	NAND3X1 NAND3X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_14749_), .B(_14783_), .C(_14717_), .Y(_14794_) );
	NOR2X1 NOR2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_14662_), .B(_14706_), .Y(_14805_) );
	AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_14706_), .B(_14662_), .Y(_14815_) );
	OAI21X1 OAI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_14805_), .B(_14815_), .C(_14772_), .Y(_14826_) );
	NAND3X1 NAND3X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_13808_), .B(_14794_), .C(_14826_), .Y(_14837_) );
	NAND3X1 NAND3X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_14749_), .B(_14772_), .C(_14717_), .Y(_14848_) );
	OAI21X1 OAI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_14805_), .B(_14815_), .C(_14783_), .Y(_14859_) );
	NAND3X1 NAND3X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_13819_), .B(_14848_), .C(_14859_), .Y(_14870_) );
	AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_14837_), .B(_14870_), .Y(_14881_) );
	AOI21X1 AOI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_14115_), .B(_14071_), .C(_13994_), .Y(_14892_) );
	OAI21X1 OAI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_14192_), .B(_14892_), .C(_14126_), .Y(_14903_) );
	NOR2X1 NOR2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_13436__bF_buf1), .Y(_14914_) );
	NAND2X1 NAND2X1_2438 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf5), .B(aOperand_frameOut_5_bF_buf1), .Y(_14925_) );
	OAI21X1 OAI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf0), .B(_12780_), .C(_13939_), .Y(_14936_) );
	OAI21X1 OAI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_14760_), .B(_14925_), .C(_14936_), .Y(_14947_) );
	XNOR2X1 XNOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_14947_), .B(_14914_), .Y(_14958_) );
	AOI21X1 AOI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_14060_), .B(_14005_), .C(_14037_), .Y(_14969_) );
	INVX1 INVX1_1673 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .Y(_14980_) );
	NAND2X1 NAND2X1_2439 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf3), .B(aOperand_frameOut_6_bF_buf3), .Y(_14991_) );
	INVX1 INVX1_1674 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .Y(_15002_) );
	NAND2X1 NAND2X1_2440 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_8_bF_buf0), .Y(_15013_) );
	OR2X2 OR2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_14093_), .B(_15013_), .Y(_15024_) );
	INVX8 INVX8_62 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf4), .Y(_15035_) );
	OAI21X1 OAI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf3), .B(_15035_), .C(_14093_), .Y(_15046_) );
	NAND3X1 NAND3X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_15002_), .B(_15046_), .C(_15024_), .Y(_15057_) );
	NOR2X1 NOR2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_14093_), .B(_15013_), .Y(_15068_) );
	AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_14093_), .B(_15013_), .Y(_15079_) );
	OAI21X1 OAI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_15068_), .B(_15079_), .C(_14991_), .Y(_15090_) );
	NAND3X1 NAND3X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_15057_), .B(_15090_), .C(_14980_), .Y(_15101_) );
	NOR3X1 NOR3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .B(_15068_), .C(_15079_), .Y(_15112_) );
	AOI21X1 AOI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_15024_), .B(_15046_), .C(_15002_), .Y(_15122_) );
	OAI21X1 OAI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_15122_), .B(_15112_), .C(_14969_), .Y(_15133_) );
	NAND3X1 NAND3X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_14958_), .B(_15133_), .C(_15101_), .Y(_15144_) );
	XOR2X1 XOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_14947_), .B(_14914_), .Y(_15155_) );
	OAI21X1 OAI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_15122_), .B(_15112_), .C(_14980_), .Y(_15166_) );
	NAND3X1 NAND3X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .B(_15090_), .C(_15057_), .Y(_15177_) );
	NAND3X1 NAND3X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_15155_), .C(_15166_), .Y(_15188_) );
	NAND3X1 NAND3X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_15144_), .B(_15188_), .C(_14903_), .Y(_15199_) );
	INVX1 INVX1_1675 ( .gnd(gnd), .vdd(vdd), .A(_14126_), .Y(_15210_) );
	AOI21X1 AOI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_13972_), .B(_14170_), .C(_15210_), .Y(_15221_) );
	AOI21X1 AOI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_15166_), .B(_15177_), .C(_15155_), .Y(_15232_) );
	AOI21X1 AOI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_15101_), .B(_15133_), .C(_14958_), .Y(_15243_) );
	OAI21X1 OAI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_15232_), .B(_15243_), .C(_15221_), .Y(_15264_) );
	NAND3X1 NAND3X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_15199_), .B(_14881_), .C(_15264_), .Y(_15265_) );
	NAND2X1 NAND2X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_14837_), .B(_14870_), .Y(_15276_) );
	OAI21X1 OAI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_15232_), .B(_15243_), .C(_14903_), .Y(_15287_) );
	NAND3X1 NAND3X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_15144_), .B(_15188_), .C(_15221_), .Y(_15298_) );
	NAND3X1 NAND3X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_15276_), .B(_15287_), .C(_15298_), .Y(_15309_) );
	NAND3X1 NAND3X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_15265_), .B(_15309_), .C(_14651_), .Y(_15320_) );
	NAND2X1 NAND2X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_14225_), .B(_14181_), .Y(_15331_) );
	NOR2X1 NOR2X1_800 ( .gnd(gnd), .vdd(vdd), .A(_14257_), .B(_15331_), .Y(_15342_) );
	AOI21X1 AOI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_13896_), .B(_14290_), .C(_15342_), .Y(_15353_) );
	AOI21X1 AOI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_15298_), .B(_15287_), .C(_15276_), .Y(_15364_) );
	AOI21X1 AOI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_15264_), .B(_15199_), .C(_14881_), .Y(_15375_) );
	OAI21X1 OAI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_15375_), .B(_15364_), .C(_15353_), .Y(_15386_) );
	NAND3X1 NAND3X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_14629_), .B(_15320_), .C(_15386_), .Y(_15397_) );
	OAI21X1 OAI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_15375_), .B(_15364_), .C(_14651_), .Y(_15408_) );
	NAND3X1 NAND3X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_15265_), .B(_15309_), .C(_15353_), .Y(_15419_) );
	NAND3X1 NAND3X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_15408_), .C(_15419_), .Y(_15430_) );
	NAND3X1 NAND3X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_15397_), .B(_15430_), .C(_14607_), .Y(_15441_) );
	INVX1 INVX1_1676 ( .gnd(gnd), .vdd(vdd), .A(_14345_), .Y(_15451_) );
	AOI21X1 AOI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_14389_), .C(_15451_), .Y(_15462_) );
	AOI21X1 AOI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_15419_), .B(_15408_), .C(_14618_), .Y(_15473_) );
	AOI21X1 AOI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_15386_), .B(_15320_), .C(_14629_), .Y(_15484_) );
	OAI21X1 OAI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_15484_), .B(_15473_), .C(_15462_), .Y(_15495_) );
	NAND3X1 NAND3X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .B(_15495_), .C(_14585_), .Y(_15506_) );
	OAI21X1 OAI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_15484_), .B(_15473_), .C(_14607_), .Y(_15517_) );
	NAND3X1 NAND3X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_15397_), .B(_15430_), .C(_15462_), .Y(_15528_) );
	NAND3X1 NAND3X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_14552_), .B(_15528_), .C(_15517_), .Y(_15539_) );
	NAND3X1 NAND3X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_14574_), .B(_15506_), .C(_15539_), .Y(_15560_) );
	NAND2X1 NAND2X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_13677_), .B(_13655_), .Y(_15571_) );
	AOI21X1 AOI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_14444_), .B(_14498_), .C(_15571_), .Y(_15572_) );
	NAND3X1 NAND3X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .B(_14552_), .C(_15495_), .Y(_15583_) );
	NAND3X1 NAND3X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_15528_), .B(_14585_), .C(_15517_), .Y(_15594_) );
	NAND3X1 NAND3X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_15583_), .B(_15594_), .C(_15572_), .Y(_15605_) );
	AOI21X1 AOI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_15605_), .B(_15560_), .C(_14541_), .Y(_15616_) );
	INVX1 INVX1_1677 ( .gnd(gnd), .vdd(vdd), .A(_15616_), .Y(_15627_) );
	NAND3X1 NAND3X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_15560_), .B(_15605_), .C(_14541_), .Y(_15638_) );
	AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_15627_), .B(_15638_), .Y(mulOut_8_) );
	NAND3X1 NAND3X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_15506_), .B(_15539_), .C(_15572_), .Y(_15659_) );
	INVX1 INVX1_1678 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .Y(_15670_) );
	AOI21X1 AOI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_15309_), .B(_15265_), .C(_14651_), .Y(_15681_) );
	OAI21X1 OAI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_15681_), .C(_15320_), .Y(_15692_) );
	AOI21X1 AOI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_15144_), .B(_15188_), .C(_14903_), .Y(_15703_) );
	OAI21X1 OAI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_15276_), .B(_15703_), .C(_15199_), .Y(_15714_) );
	AOI21X1 AOI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_15057_), .B(_15090_), .C(_14980_), .Y(_15725_) );
	OAI21X1 OAI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_15155_), .B(_15725_), .C(_15101_), .Y(_15736_) );
	OAI21X1 OAI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .B(_15079_), .C(_15024_), .Y(_15747_) );
	NAND2X1 NAND2X1_2444 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf2), .B(aOperand_frameOut_7_bF_buf3), .Y(_15758_) );
	INVX1 INVX1_1679 ( .gnd(gnd), .vdd(vdd), .A(_15758_), .Y(_15769_) );
	AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf4), .B(aOperand_frameOut_8_bF_buf3), .Y(_15779_) );
	AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_9_bF_buf4), .Y(_15790_) );
	NAND2X1 NAND2X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_15779_), .B(_15790_), .Y(_15801_) );
	INVX8 INVX8_63 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf3), .Y(_15812_) );
	OAI22X1 OAI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf2), .B(_15812__bF_buf3), .C(_11776__bF_buf1), .D(_15035_), .Y(_15823_) );
	NAND3X1 NAND3X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_15769_), .B(_15823_), .C(_15801_), .Y(_15834_) );
	OAI21X1 OAI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf0), .B(_15035_), .C(_15790_), .Y(_15845_) );
	OAI21X1 OAI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf1), .B(_15812__bF_buf2), .C(_15779_), .Y(_15856_) );
	NAND3X1 NAND3X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_15758_), .B(_15845_), .C(_15856_), .Y(_15867_) );
	NAND3X1 NAND3X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .B(_15867_), .C(_15747_), .Y(_15878_) );
	AOI21X1 AOI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_15046_), .B(_15002_), .C(_15068_), .Y(_15889_) );
	AOI21X1 AOI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_15845_), .B(_15856_), .C(_15758_), .Y(_15900_) );
	AOI21X1 AOI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_15801_), .B(_15823_), .C(_15769_), .Y(_15911_) );
	OAI21X1 OAI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_15911_), .B(_15900_), .C(_15889_), .Y(_15922_) );
	NAND2X1 NAND2X1_2446 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf1), .B(adder_bOperand_5_bF_buf1), .Y(_15933_) );
	INVX1 INVX1_1680 ( .gnd(gnd), .vdd(vdd), .A(_15933_), .Y(_15944_) );
	NAND2X1 NAND2X1_2447 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .B(aOperand_frameOut_5_bF_buf0), .Y(_15955_) );
	NAND2X1 NAND2X1_2448 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .B(aOperand_frameOut_6_bF_buf2), .Y(_15966_) );
	OAI21X1 OAI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf3), .B(_13294__bF_buf2), .C(_14925_), .Y(_15977_) );
	OAI21X1 OAI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15966_), .C(_15977_), .Y(_15988_) );
	XNOR2X1 XNOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_15988_), .B(_15944_), .Y(_15999_) );
	NAND3X1 NAND3X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_15922_), .B(_15878_), .C(_15999_), .Y(_16010_) );
	OAI21X1 OAI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_15911_), .B(_15900_), .C(_15747_), .Y(_16021_) );
	NAND3X1 NAND3X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .B(_15889_), .C(_15867_), .Y(_16032_) );
	XNOR2X1 XNOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_15988_), .B(_15933_), .Y(_16043_) );
	NAND3X1 NAND3X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_16021_), .B(_16032_), .C(_16043_), .Y(_16054_) );
	NAND3X1 NAND3X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_16010_), .B(_16054_), .C(_15736_), .Y(_16065_) );
	NAND2X1 NAND2X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_15090_), .B(_15057_), .Y(_16075_) );
	NOR2X1 NOR2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .B(_16075_), .Y(_16096_) );
	AOI21X1 AOI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_15133_), .B(_14958_), .C(_16096_), .Y(_16097_) );
	AOI21X1 AOI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_16021_), .B(_16032_), .C(_16043_), .Y(_16108_) );
	AOI21X1 AOI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_15922_), .B(_15878_), .C(_15999_), .Y(_16119_) );
	OAI21X1 OAI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_16108_), .B(_16119_), .C(_16097_), .Y(_16130_) );
	NAND2X1 NAND2X1_2450 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf4), .B(adder_bOperand_6_bF_buf5), .Y(_16141_) );
	NOR2X1 NOR2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_13797_), .B(_16141_), .Y(_16152_) );
	NOR2X1 NOR2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_16152_), .B(_14805_), .Y(_16163_) );
	NAND2X1 NAND2X1_2451 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf5), .B(adder_bOperand_8_bF_buf3), .Y(_16174_) );
	NAND2X1 NAND2X1_2452 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf0), .B(adder_bOperand_7_bF_buf0), .Y(_16185_) );
	OAI21X1 OAI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_14684__bF_buf2), .C(_14673_), .Y(_16196_) );
	OAI21X1 OAI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_16141_), .B(_16185_), .C(_16196_), .Y(_16207_) );
	OR2X2 OR2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_16207_), .B(_16174_), .Y(_16218_) );
	OAI21X1 OAI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_14728__bF_buf2), .C(_16207_), .Y(_16229_) );
	NOR2X1 NOR2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_13939_), .B(_15955_), .Y(_16240_) );
	AOI21X1 AOI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .B(_14914_), .C(_16240_), .Y(_16251_) );
	INVX1 INVX1_1681 ( .gnd(gnd), .vdd(vdd), .A(_16251_), .Y(_16262_) );
	NAND3X1 NAND3X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_16229_), .B(_16262_), .C(_16218_), .Y(_16273_) );
	NOR2X1 NOR2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_16174_), .B(_16207_), .Y(_16284_) );
	AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_16207_), .B(_16174_), .Y(_16295_) );
	OAI21X1 OAI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_16284_), .B(_16295_), .C(_16251_), .Y(_16306_) );
	NAND3X1 NAND3X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_16273_), .C(_16306_), .Y(_16317_) );
	OAI21X1 OAI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_13797_), .B(_16141_), .C(_14717_), .Y(_16328_) );
	NAND3X1 NAND3X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_16229_), .B(_16251_), .C(_16218_), .Y(_16339_) );
	OAI21X1 OAI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_16284_), .B(_16295_), .C(_16262_), .Y(_16350_) );
	NAND3X1 NAND3X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_16328_), .B(_16339_), .C(_16350_), .Y(_16360_) );
	NAND2X1 NAND2X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_16317_), .B(_16360_), .Y(_16371_) );
	NAND3X1 NAND3X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_16065_), .B(_16371_), .C(_16130_), .Y(_16382_) );
	OAI21X1 OAI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_16108_), .B(_16119_), .C(_15736_), .Y(_16403_) );
	NAND3X1 NAND3X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_16010_), .B(_16054_), .C(_16097_), .Y(_16414_) );
	NAND3X1 NAND3X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_16328_), .B(_16273_), .C(_16306_), .Y(_16415_) );
	NAND3X1 NAND3X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_16339_), .C(_16350_), .Y(_16426_) );
	NAND2X1 NAND2X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_16426_), .B(_16415_), .Y(_16437_) );
	NAND3X1 NAND3X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_16403_), .B(_16437_), .C(_16414_), .Y(_16448_) );
	NAND3X1 NAND3X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_16448_), .B(_16382_), .C(_15714_), .Y(_16459_) );
	INVX1 INVX1_1682 ( .gnd(gnd), .vdd(vdd), .A(_15714_), .Y(_16470_) );
	AOI21X1 AOI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_16414_), .B(_16403_), .C(_16437_), .Y(_16481_) );
	AOI21X1 AOI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_16130_), .B(_16065_), .C(_16371_), .Y(_16492_) );
	OAI21X1 OAI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_16481_), .B(_16492_), .C(_16470_), .Y(_16503_) );
	NAND2X1 NAND2X1_2455 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf3), .B(adder_bOperand_9_bF_buf1), .Y(_16514_) );
	INVX1 INVX1_1683 ( .gnd(gnd), .vdd(vdd), .A(_16514_), .Y(_16525_) );
	NAND2X1 NAND2X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_14794_), .B(_14837_), .Y(_16536_) );
	XNOR2X1 XNOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_16536_), .B(_16525_), .Y(_16547_) );
	INVX1 INVX1_1684 ( .gnd(gnd), .vdd(vdd), .A(_16547_), .Y(_16558_) );
	NAND3X1 NAND3X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_16459_), .B(_16558_), .C(_16503_), .Y(_16569_) );
	INVX1 INVX1_1685 ( .gnd(gnd), .vdd(vdd), .A(_16459_), .Y(_16580_) );
	AOI21X1 AOI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_16382_), .B(_16448_), .C(_15714_), .Y(_16591_) );
	OAI21X1 OAI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_16591_), .B(_16580_), .C(_16547_), .Y(_16602_) );
	NAND3X1 NAND3X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_15692_), .B(_16569_), .C(_16602_), .Y(_16613_) );
	INVX1 INVX1_1686 ( .gnd(gnd), .vdd(vdd), .A(_15692_), .Y(_16624_) );
	NOR3X1 NOR3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_16591_), .B(_16547_), .C(_16580_), .Y(_16635_) );
	AOI21X1 AOI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_16503_), .B(_16459_), .C(_16558_), .Y(_16645_) );
	OAI21X1 OAI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_16645_), .B(_16635_), .C(_16624_), .Y(_16656_) );
	NAND3X1 NAND3X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_16613_), .B(_16656_), .C(_15670_), .Y(_16667_) );
	OAI21X1 OAI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_16645_), .B(_16635_), .C(_15692_), .Y(_16678_) );
	NAND3X1 NAND3X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_16569_), .B(_16602_), .C(_16624_), .Y(_16689_) );
	NAND3X1 NAND3X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .B(_16678_), .C(_16689_), .Y(_16700_) );
	NAND2X1 NAND2X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_16700_), .B(_16667_), .Y(_16711_) );
	NAND3X1 NAND3X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_15506_), .B(_16711_), .C(_15659_), .Y(_16722_) );
	AOI21X1 AOI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_16689_), .B(_16678_), .C(_15441_), .Y(_16733_) );
	NOR2X1 NOR2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_15484_), .B(_15473_), .Y(_16744_) );
	AOI22X1 AOI22X1_271 ( .gnd(gnd), .vdd(vdd), .A(_16744_), .B(_14607_), .C(_16613_), .D(_16656_), .Y(_16755_) );
	NOR2X1 NOR2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_16755_), .B(_16733_), .Y(_16766_) );
	AOI21X1 AOI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_15495_), .B(_15441_), .C(_14585_), .Y(_16777_) );
	OAI21X1 OAI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_14574_), .B(_16777_), .C(_15506_), .Y(_16788_) );
	NAND2X1 NAND2X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_16788_), .B(_16766_), .Y(_16799_) );
	NAND3X1 NAND3X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_16722_), .B(_16799_), .C(_15616_), .Y(_16810_) );
	INVX1 INVX1_1687 ( .gnd(gnd), .vdd(vdd), .A(_16810_), .Y(_16821_) );
	INVX1 INVX1_1688 ( .gnd(gnd), .vdd(vdd), .A(_16613_), .Y(_16832_) );
	NAND2X1 NAND2X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_16525_), .B(_16536_), .Y(_16843_) );
	INVX1 INVX1_1689 ( .gnd(gnd), .vdd(vdd), .A(_16843_), .Y(_16854_) );
	OAI21X1 OAI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_16547_), .B(_16591_), .C(_16459_), .Y(_16865_) );
	NAND2X1 NAND2X1_2460 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf4), .B(adder_bOperand_10_bF_buf4), .Y(_16876_) );
	INVX4 INVX4_13 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf3), .Y(_16887_) );
	NAND2X1 NAND2X1_2461 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf3), .B(adder_bOperand_9_bF_buf0), .Y(_16895_) );
	OAI21X1 OAI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf1), .B(_16887_), .C(_16895_), .Y(_16896_) );
	OAI21X1 OAI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_16514_), .B(_16876_), .C(_16896_), .Y(_16897_) );
	NAND2X1 NAND2X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_16273_), .B(_16415_), .Y(_16898_) );
	XNOR2X1 XNOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_16898_), .B(_16897_), .Y(_16899_) );
	AOI21X1 AOI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_16010_), .B(_16054_), .C(_15736_), .Y(_16900_) );
	OAI21X1 OAI21X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_16900_), .B(_16437_), .C(_16065_), .Y(_16901_) );
	INVX1 INVX1_1690 ( .gnd(gnd), .vdd(vdd), .A(_16141_), .Y(_16902_) );
	INVX1 INVX1_1691 ( .gnd(gnd), .vdd(vdd), .A(_16185_), .Y(_16903_) );
	AOI21X1 AOI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_16902_), .B(_16903_), .C(_16284_), .Y(_16904_) );
	NAND2X1 NAND2X1_2463 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf3), .B(adder_bOperand_8_bF_buf2), .Y(_16905_) );
	NAND2X1 NAND2X1_2464 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf4), .B(adder_bOperand_6_bF_buf4), .Y(_16906_) );
	NAND2X1 NAND2X1_2465 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf0), .B(adder_bOperand_7_bF_buf5), .Y(_16907_) );
	OAI21X1 OAI21X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf3), .B(_14684__bF_buf1), .C(_16185_), .Y(_16908_) );
	OAI21X1 OAI21X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_16906_), .B(_16907_), .C(_16908_), .Y(_16909_) );
	OR2X2 OR2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_16909_), .B(_16905_), .Y(_16910_) );
	OAI21X1 OAI21X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf3), .B(_14728__bF_buf1), .C(_16909_), .Y(_16911_) );
	NAND2X1 NAND2X1_2466 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf3), .B(aOperand_frameOut_6_bF_buf1), .Y(_16912_) );
	NOR2X1 NOR2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_14925_), .B(_16912_), .Y(_16913_) );
	AOI21X1 AOI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_15977_), .B(_15944_), .C(_16913_), .Y(_16914_) );
	INVX1 INVX1_1692 ( .gnd(gnd), .vdd(vdd), .A(_16914_), .Y(_16915_) );
	NAND3X1 NAND3X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_16911_), .B(_16915_), .C(_16910_), .Y(_16916_) );
	NOR2X1 NOR2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_16905_), .B(_16909_), .Y(_16917_) );
	AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_16909_), .B(_16905_), .Y(_16918_) );
	OAI21X1 OAI21X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_16917_), .B(_16918_), .C(_16914_), .Y(_16919_) );
	NAND3X1 NAND3X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_16904_), .B(_16916_), .C(_16919_), .Y(_16920_) );
	OAI21X1 OAI21X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_16141_), .B(_16185_), .C(_16218_), .Y(_16921_) );
	NAND3X1 NAND3X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_16911_), .B(_16914_), .C(_16910_), .Y(_16922_) );
	OAI21X1 OAI21X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_16917_), .B(_16918_), .C(_16915_), .Y(_16923_) );
	NAND3X1 NAND3X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_16921_), .B(_16922_), .C(_16923_), .Y(_16924_) );
	NAND2X1 NAND2X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_16920_), .B(_16924_), .Y(_16925_) );
	AOI21X1 AOI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_15867_), .B(_15834_), .C(_15747_), .Y(_16926_) );
	OAI21X1 OAI21X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_16926_), .B(_16043_), .C(_15878_), .Y(_16927_) );
	NOR2X1 NOR2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_13436__bF_buf0), .Y(_16928_) );
	NAND2X1 NAND2X1_2468 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf3), .B(aOperand_frameOut_7_bF_buf2), .Y(_16929_) );
	OAI21X1 OAI21X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf2), .B(_14049_), .C(_15966_), .Y(_16930_) );
	OAI21X1 OAI21X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_16912_), .B(_16929_), .C(_16930_), .Y(_16931_) );
	XNOR2X1 XNOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_16931_), .B(_16928_), .Y(_16932_) );
	NOR2X1 NOR2X1_811 ( .gnd(gnd), .vdd(vdd), .A(_15779_), .B(_15790_), .Y(_16933_) );
	OAI21X1 OAI21X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_15758_), .B(_16933_), .C(_15801_), .Y(_16934_) );
	NAND2X1 NAND2X1_2469 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf1), .B(aOperand_frameOut_8_bF_buf2), .Y(_16935_) );
	INVX1 INVX1_1693 ( .gnd(gnd), .vdd(vdd), .A(_16935_), .Y(_16936_) );
	AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf3), .B(aOperand_frameOut_9_bF_buf2), .Y(_16937_) );
	AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_10_bF_buf0), .Y(_16938_) );
	NAND2X1 NAND2X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_16937_), .B(_16938_), .Y(_16939_) );
	INVX8 INVX8_64 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf4), .Y(_16940_) );
	OAI22X1 OAI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf0), .B(_16940_), .C(_11776__bF_buf3), .D(_15812__bF_buf1), .Y(_16941_) );
	NAND3X1 NAND3X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_16936_), .B(_16941_), .C(_16939_), .Y(_16942_) );
	AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_16937_), .B(_16938_), .Y(_16943_) );
	NOR2X1 NOR2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_16937_), .B(_16938_), .Y(_16944_) );
	OAI21X1 OAI21X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_16944_), .B(_16943_), .C(_16935_), .Y(_16945_) );
	NAND3X1 NAND3X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_16942_), .B(_16934_), .C(_16945_), .Y(_16946_) );
	INVX1 INVX1_1694 ( .gnd(gnd), .vdd(vdd), .A(_15013_), .Y(_16947_) );
	AOI22X1 AOI22X1_272 ( .gnd(gnd), .vdd(vdd), .A(_16947_), .B(_16937_), .C(_15769_), .D(_15823_), .Y(_16948_) );
	OAI21X1 OAI21X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf2), .B(_15812__bF_buf0), .C(_16938_), .Y(_16949_) );
	OAI21X1 OAI21X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf4), .B(_16940_), .C(_16937_), .Y(_16950_) );
	AOI21X1 AOI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_16949_), .B(_16950_), .C(_16935_), .Y(_16951_) );
	AOI21X1 AOI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_16939_), .B(_16941_), .C(_16936_), .Y(_16952_) );
	OAI21X1 OAI21X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_16952_), .B(_16951_), .C(_16948_), .Y(_16953_) );
	NAND3X1 NAND3X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_16953_), .B(_16946_), .C(_16932_), .Y(_16954_) );
	XOR2X1 XOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_16931_), .B(_16928_), .Y(_16955_) );
	OAI21X1 OAI21X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_16952_), .B(_16951_), .C(_16934_), .Y(_16956_) );
	NAND3X1 NAND3X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_16948_), .B(_16942_), .C(_16945_), .Y(_16957_) );
	NAND3X1 NAND3X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_16956_), .B(_16957_), .C(_16955_), .Y(_16958_) );
	NAND3X1 NAND3X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_16954_), .B(_16958_), .C(_16927_), .Y(_16959_) );
	INVX1 INVX1_1695 ( .gnd(gnd), .vdd(vdd), .A(_15878_), .Y(_16960_) );
	AOI21X1 AOI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_15999_), .B(_15922_), .C(_16960_), .Y(_16961_) );
	AOI21X1 AOI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_16957_), .B(_16956_), .C(_16955_), .Y(_16962_) );
	AOI21X1 AOI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_16946_), .B(_16953_), .C(_16932_), .Y(_16963_) );
	OAI21X1 OAI21X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_16962_), .B(_16963_), .C(_16961_), .Y(_16964_) );
	NAND3X1 NAND3X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_16959_), .B(_16964_), .C(_16925_), .Y(_16965_) );
	NAND3X1 NAND3X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_16921_), .B(_16916_), .C(_16919_), .Y(_16966_) );
	NAND3X1 NAND3X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_16904_), .B(_16922_), .C(_16923_), .Y(_16967_) );
	NAND2X1 NAND2X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_16967_), .B(_16966_), .Y(_16968_) );
	OAI21X1 OAI21X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_16962_), .B(_16963_), .C(_16927_), .Y(_16969_) );
	NAND3X1 NAND3X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_16954_), .B(_16958_), .C(_16961_), .Y(_16970_) );
	NAND3X1 NAND3X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_16970_), .B(_16969_), .C(_16968_), .Y(_16971_) );
	NAND3X1 NAND3X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_16965_), .B(_16971_), .C(_16901_), .Y(_16972_) );
	NAND2X1 NAND2X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_16010_), .B(_16054_), .Y(_16973_) );
	NOR2X1 NOR2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_16097_), .B(_16973_), .Y(_16974_) );
	AOI21X1 AOI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_16130_), .B(_16371_), .C(_16974_), .Y(_16975_) );
	AOI21X1 AOI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_16969_), .B(_16970_), .C(_16968_), .Y(_16976_) );
	AOI21X1 AOI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_16964_), .B(_16959_), .C(_16925_), .Y(_16977_) );
	OAI21X1 OAI21X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_16976_), .B(_16977_), .C(_16975_), .Y(_16978_) );
	NAND3X1 NAND3X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_16899_), .B(_16972_), .C(_16978_), .Y(_16979_) );
	INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(_16897_), .Y(_16980_) );
	XNOR2X1 XNOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_16898_), .B(_16980_), .Y(_16981_) );
	OAI21X1 OAI21X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_16976_), .B(_16977_), .C(_16901_), .Y(_16982_) );
	NAND3X1 NAND3X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_16965_), .B(_16971_), .C(_16975_), .Y(_16983_) );
	NAND3X1 NAND3X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_16981_), .B(_16982_), .C(_16983_), .Y(_16984_) );
	NAND3X1 NAND3X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_16979_), .B(_16865_), .C(_16984_), .Y(_16985_) );
	AOI21X1 AOI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_16503_), .B(_16558_), .C(_16580_), .Y(_16986_) );
	AOI21X1 AOI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_16983_), .B(_16982_), .C(_16981_), .Y(_16987_) );
	AOI21X1 AOI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_16978_), .B(_16972_), .C(_16899_), .Y(_16988_) );
	OAI21X1 OAI21X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_16988_), .B(_16987_), .C(_16986_), .Y(_16989_) );
	NAND3X1 NAND3X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_16854_), .B(_16985_), .C(_16989_), .Y(_16990_) );
	OAI21X1 OAI21X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_16988_), .B(_16987_), .C(_16865_), .Y(_16991_) );
	NAND3X1 NAND3X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_16979_), .B(_16984_), .C(_16986_), .Y(_16992_) );
	NAND3X1 NAND3X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_16843_), .B(_16991_), .C(_16992_), .Y(_16993_) );
	NAND3X1 NAND3X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_16832_), .B(_16990_), .C(_16993_), .Y(_16994_) );
	NAND3X1 NAND3X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_16843_), .B(_16985_), .C(_16989_), .Y(_16995_) );
	NAND3X1 NAND3X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_16854_), .B(_16991_), .C(_16992_), .Y(_16996_) );
	NAND3X1 NAND3X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_16613_), .B(_16995_), .C(_16996_), .Y(_16997_) );
	NAND2X1 NAND2X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_16997_), .B(_16994_), .Y(_16998_) );
	AOI21X1 AOI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_15517_), .B(_15528_), .C(_14552_), .Y(_16999_) );
	AOI21X1 AOI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_16999_), .B(_16700_), .C(_16733_), .Y(_17000_) );
	NAND2X1 NAND2X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_17000_), .B(_16998_), .Y(_17001_) );
	NAND3X1 NAND3X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_16613_), .B(_16990_), .C(_16993_), .Y(_17002_) );
	NAND3X1 NAND3X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_16832_), .B(_16995_), .C(_16996_), .Y(_17003_) );
	NAND2X1 NAND2X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_17002_), .B(_17003_), .Y(_17004_) );
	OAI21X1 OAI21X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_15506_), .B(_16755_), .C(_16667_), .Y(_17005_) );
	NAND2X1 NAND2X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_17005_), .B(_17004_), .Y(_17006_) );
	NOR2X1 NOR2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_16711_), .B(_15659_), .Y(_17007_) );
	NAND3X1 NAND3X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_17007_), .B(_17006_), .C(_17001_), .Y(_17008_) );
	INVX1 INVX1_1696 ( .gnd(gnd), .vdd(vdd), .A(_15659_), .Y(_17009_) );
	AOI22X1 AOI22X1_273 ( .gnd(gnd), .vdd(vdd), .A(_17009_), .B(_16766_), .C(_17006_), .D(_17001_), .Y(_17010_) );
	INVX1 INVX1_1697 ( .gnd(gnd), .vdd(vdd), .A(_17010_), .Y(_17011_) );
	NAND2X1 NAND2X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_17008_), .B(_17011_), .Y(_17012_) );
	XNOR2X1 XNOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_17012_), .B(_16821_), .Y(mulOut_10_) );
	NAND3X1 NAND3X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_16999_), .B(_16766_), .C(_17004_), .Y(_17013_) );
	NAND3X1 NAND3X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_16733_), .B(_16997_), .C(_16994_), .Y(_17014_) );
	AOI21X1 AOI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_16996_), .B(_16995_), .C(_16613_), .Y(_17015_) );
	AOI21X1 AOI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_16984_), .B(_16979_), .C(_16865_), .Y(_17016_) );
	OAI21X1 OAI21X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_16843_), .B(_17016_), .C(_16985_), .Y(_17017_) );
	NAND2X1 NAND2X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_16980_), .B(_16898_), .Y(_17018_) );
	INVX1 INVX1_1698 ( .gnd(gnd), .vdd(vdd), .A(_17018_), .Y(_17019_) );
	AOI21X1 AOI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_16971_), .B(_16965_), .C(_16901_), .Y(_17020_) );
	OAI21X1 OAI21X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_16981_), .B(_17020_), .C(_16972_), .Y(_17021_) );
	INVX8 INVX8_65 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf3), .Y(_17022_) );
	NOR2X1 NOR2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf0), .B(_17022__bF_buf3), .Y(_17023_) );
	NAND2X1 NAND2X1_2479 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf2), .B(adder_bOperand_10_bF_buf2), .Y(_17024_) );
	INVX8 INVX8_66 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf4), .Y(_17025_) );
	OAI21X1 OAI21X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf2), .B(_17025__bF_buf3), .C(_16876_), .Y(_17026_) );
	OAI21X1 OAI21X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_16895_), .B(_17024_), .C(_17026_), .Y(_17027_) );
	XOR2X1 XOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_17027_), .B(_17023_), .Y(_17028_) );
	OAI21X1 OAI21X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_16514_), .B(_16876_), .C(_17028_), .Y(_17029_) );
	NOR2X1 NOR2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_16514_), .B(_16876_), .Y(_17030_) );
	INVX1 INVX1_1699 ( .gnd(gnd), .vdd(vdd), .A(_17030_), .Y(_17031_) );
	NOR2X1 NOR2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_17031_), .B(_17028_), .Y(_17032_) );
	INVX1 INVX1_1700 ( .gnd(gnd), .vdd(vdd), .A(_17032_), .Y(_17033_) );
	NAND2X1 NAND2X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_17029_), .B(_17033_), .Y(_17034_) );
	AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_16966_), .B(_16916_), .Y(_17035_) );
	XOR2X1 XOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_17035_), .B(_17034_), .Y(_17036_) );
	AOI21X1 AOI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_16958_), .B(_16954_), .C(_16927_), .Y(_17037_) );
	OAI21X1 OAI21X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_17037_), .B(_16968_), .C(_16959_), .Y(_17038_) );
	NAND2X1 NAND2X1_2481 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf4), .B(adder_bOperand_6_bF_buf3), .Y(_17039_) );
	INVX1 INVX1_1701 ( .gnd(gnd), .vdd(vdd), .A(_17039_), .Y(_17040_) );
	AOI21X1 AOI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_16903_), .B(_17040_), .C(_16917_), .Y(_17041_) );
	NAND2X1 NAND2X1_2482 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf3), .B(adder_bOperand_8_bF_buf1), .Y(_17042_) );
	NAND2X1 NAND2X1_2483 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf4), .B(adder_bOperand_7_bF_buf4), .Y(_17043_) );
	OAI21X1 OAI21X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_14684__bF_buf0), .C(_16907_), .Y(_17044_) );
	OAI21X1 OAI21X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_17039_), .B(_17043_), .C(_17044_), .Y(_17045_) );
	OR2X2 OR2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_17045_), .B(_17042_), .Y(_17046_) );
	OAI21X1 OAI21X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_14728__bF_buf0), .C(_17045_), .Y(_17047_) );
	NAND2X1 NAND2X1_2484 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf2), .B(aOperand_frameOut_7_bF_buf1), .Y(_17048_) );
	NOR2X1 NOR2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_15966_), .B(_17048_), .Y(_17049_) );
	AOI21X1 AOI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_16930_), .B(_16928_), .C(_17049_), .Y(_17050_) );
	INVX1 INVX1_1702 ( .gnd(gnd), .vdd(vdd), .A(_17050_), .Y(_17051_) );
	NAND3X1 NAND3X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_17047_), .B(_17051_), .C(_17046_), .Y(_17052_) );
	NOR2X1 NOR2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_17042_), .B(_17045_), .Y(_17053_) );
	AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_17045_), .B(_17042_), .Y(_17054_) );
	OAI21X1 OAI21X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_17053_), .B(_17054_), .C(_17050_), .Y(_17055_) );
	NAND3X1 NAND3X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_17041_), .B(_17052_), .C(_17055_), .Y(_17056_) );
	OAI21X1 OAI21X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_16906_), .B(_16907_), .C(_16910_), .Y(_17057_) );
	NAND3X1 NAND3X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_17047_), .B(_17050_), .C(_17046_), .Y(_17058_) );
	OAI21X1 OAI21X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_17053_), .B(_17054_), .C(_17051_), .Y(_17059_) );
	NAND3X1 NAND3X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_17057_), .B(_17058_), .C(_17059_), .Y(_17060_) );
	NAND2X1 NAND2X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_17056_), .B(_17060_), .Y(_17061_) );
	AOI21X1 AOI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_16945_), .B(_16942_), .C(_16934_), .Y(_17062_) );
	OAI21X1 OAI21X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_16955_), .B(_17062_), .C(_16946_), .Y(_17063_) );
	NOR2X1 NOR2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf3), .B(_13294__bF_buf1), .Y(_17064_) );
	NAND2X1 NAND2X1_2486 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf2), .B(aOperand_frameOut_8_bF_buf1), .Y(_17065_) );
	OAI21X1 OAI21X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf1), .B(_15035_), .C(_16929_), .Y(_17066_) );
	OAI21X1 OAI21X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_17048_), .B(_17065_), .C(_17066_), .Y(_17067_) );
	OR2X2 OR2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_17067_), .B(_17064_), .Y(_17068_) );
	NAND2X1 NAND2X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_17064_), .B(_17067_), .Y(_17069_) );
	NAND2X1 NAND2X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_17069_), .B(_17068_), .Y(_17070_) );
	OAI21X1 OAI21X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_16935_), .B(_16944_), .C(_16939_), .Y(_17071_) );
	NAND2X1 NAND2X1_2489 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf0), .B(aOperand_frameOut_9_bF_buf1), .Y(_17072_) );
	INVX1 INVX1_1703 ( .gnd(gnd), .vdd(vdd), .A(_17072_), .Y(_17073_) );
	NAND2X1 NAND2X1_2490 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .B(aOperand_frameOut_10_bF_buf3), .Y(_17074_) );
	NAND2X1 NAND2X1_2491 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(aOperand_frameOut_11_bF_buf2), .Y(_17075_) );
	OR2X2 OR2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_17074_), .B(_17075_), .Y(_17076_) );
	INVX8 INVX8_67 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf1), .Y(_17077_) );
	OAI21X1 OAI21X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf3), .B(_17077_), .C(_17074_), .Y(_17078_) );
	NAND3X1 NAND3X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_17073_), .B(_17078_), .C(_17076_), .Y(_17079_) );
	NOR2X1 NOR2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_17074_), .B(_17075_), .Y(_17080_) );
	AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_17074_), .B(_17075_), .Y(_17081_) );
	OAI21X1 OAI21X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_17080_), .B(_17081_), .C(_17072_), .Y(_17082_) );
	NAND3X1 NAND3X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_17079_), .B(_17082_), .C(_17071_), .Y(_17083_) );
	AOI21X1 AOI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_16941_), .B(_16936_), .C(_16943_), .Y(_17084_) );
	NOR3X1 NOR3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_17072_), .B(_17080_), .C(_17081_), .Y(_17085_) );
	AOI21X1 AOI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_17076_), .B(_17078_), .C(_17073_), .Y(_17086_) );
	OAI21X1 OAI21X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_17086_), .B(_17085_), .C(_17084_), .Y(_17087_) );
	NAND3X1 NAND3X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_17083_), .B(_17087_), .C(_17070_), .Y(_17088_) );
	XOR2X1 XOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_17067_), .B(_17064_), .Y(_17089_) );
	OAI21X1 OAI21X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_17086_), .B(_17085_), .C(_17071_), .Y(_17090_) );
	NAND3X1 NAND3X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_17079_), .B(_17082_), .C(_17084_), .Y(_17091_) );
	NAND3X1 NAND3X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_17091_), .B(_17089_), .C(_17090_), .Y(_17092_) );
	NAND3X1 NAND3X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_17092_), .B(_17088_), .C(_17063_), .Y(_17093_) );
	NOR3X1 NOR3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_16948_), .B(_16952_), .C(_16951_), .Y(_17094_) );
	AOI21X1 AOI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_16932_), .B(_16953_), .C(_17094_), .Y(_17095_) );
	AOI21X1 AOI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_17090_), .B(_17091_), .C(_17089_), .Y(_17096_) );
	AOI21X1 AOI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_17087_), .B(_17083_), .C(_17070_), .Y(_17097_) );
	OAI21X1 OAI21X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_17096_), .B(_17097_), .C(_17095_), .Y(_17098_) );
	NAND3X1 NAND3X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_17093_), .B(_17061_), .C(_17098_), .Y(_17099_) );
	NAND3X1 NAND3X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_17057_), .B(_17052_), .C(_17055_), .Y(_17100_) );
	NAND3X1 NAND3X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_17041_), .B(_17058_), .C(_17059_), .Y(_17101_) );
	NAND2X1 NAND2X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_17101_), .B(_17100_), .Y(_17102_) );
	OAI21X1 OAI21X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_17096_), .B(_17097_), .C(_17063_), .Y(_17103_) );
	NAND3X1 NAND3X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_17092_), .B(_17095_), .C(_17088_), .Y(_17104_) );
	NAND3X1 NAND3X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_17104_), .B(_17102_), .C(_17103_), .Y(_17105_) );
	NAND3X1 NAND3X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_17105_), .B(_17099_), .C(_17038_), .Y(_17106_) );
	INVX1 INVX1_1704 ( .gnd(gnd), .vdd(vdd), .A(_16959_), .Y(_17107_) );
	AOI21X1 AOI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_16925_), .B(_16964_), .C(_17107_), .Y(_17108_) );
	AOI21X1 AOI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_17103_), .B(_17104_), .C(_17102_), .Y(_17109_) );
	AOI21X1 AOI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_17098_), .B(_17093_), .C(_17061_), .Y(_17110_) );
	OAI21X1 OAI21X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_17109_), .B(_17110_), .C(_17108_), .Y(_17111_) );
	NAND3X1 NAND3X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_17106_), .B(_17036_), .C(_17111_), .Y(_17112_) );
	OR2X2 OR2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_17035_), .B(_17034_), .Y(_17113_) );
	NAND2X1 NAND2X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_17034_), .B(_17035_), .Y(_17114_) );
	NAND2X1 NAND2X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_17114_), .B(_17113_), .Y(_17115_) );
	OAI21X1 OAI21X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_17109_), .B(_17110_), .C(_17038_), .Y(_17116_) );
	NAND3X1 NAND3X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_17099_), .B(_17105_), .C(_17108_), .Y(_17117_) );
	NAND3X1 NAND3X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_17115_), .B(_17117_), .C(_17116_), .Y(_17118_) );
	NAND3X1 NAND3X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_17021_), .B(_17112_), .C(_17118_), .Y(_17119_) );
	INVX1 INVX1_1705 ( .gnd(gnd), .vdd(vdd), .A(_16972_), .Y(_17120_) );
	AOI21X1 AOI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_16899_), .B(_16978_), .C(_17120_), .Y(_17121_) );
	AOI21X1 AOI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_17116_), .B(_17117_), .C(_17115_), .Y(_17122_) );
	AOI21X1 AOI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_17111_), .B(_17106_), .C(_17036_), .Y(_17123_) );
	OAI21X1 OAI21X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_17123_), .B(_17122_), .C(_17121_), .Y(_17124_) );
	NAND3X1 NAND3X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_17019_), .B(_17119_), .C(_17124_), .Y(_17125_) );
	OAI21X1 OAI21X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_17123_), .B(_17122_), .C(_17021_), .Y(_17126_) );
	NAND3X1 NAND3X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_17112_), .B(_17118_), .C(_17121_), .Y(_17127_) );
	NAND3X1 NAND3X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_17018_), .B(_17127_), .C(_17126_), .Y(_17128_) );
	NAND3X1 NAND3X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_17017_), .B(_17125_), .C(_17128_), .Y(_17129_) );
	INVX1 INVX1_1706 ( .gnd(gnd), .vdd(vdd), .A(_16985_), .Y(_17130_) );
	AOI21X1 AOI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_16854_), .B(_16989_), .C(_17130_), .Y(_17131_) );
	AOI21X1 AOI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_17126_), .B(_17127_), .C(_17018_), .Y(_17132_) );
	AOI22X1 AOI22X1_274 ( .gnd(gnd), .vdd(vdd), .A(_16980_), .B(_16898_), .C(_17119_), .D(_17124_), .Y(_17133_) );
	OAI21X1 OAI21X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_17133_), .B(_17132_), .C(_17131_), .Y(_17134_) );
	NAND3X1 NAND3X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_17129_), .B(_17015_), .C(_17134_), .Y(_17135_) );
	OAI21X1 OAI21X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_17133_), .B(_17132_), .C(_17017_), .Y(_17136_) );
	NAND3X1 NAND3X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_17125_), .B(_17128_), .C(_17131_), .Y(_17137_) );
	NAND3X1 NAND3X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_16994_), .B(_17137_), .C(_17136_), .Y(_17138_) );
	NAND3X1 NAND3X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_17014_), .B(_17135_), .C(_17138_), .Y(_17139_) );
	AOI21X1 AOI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_17003_), .B(_17002_), .C(_16667_), .Y(_17140_) );
	NAND3X1 NAND3X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_16994_), .B(_17129_), .C(_17134_), .Y(_17141_) );
	NAND3X1 NAND3X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_17015_), .B(_17137_), .C(_17136_), .Y(_17142_) );
	NAND3X1 NAND3X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_17140_), .B(_17141_), .C(_17142_), .Y(_17143_) );
	AOI21X1 AOI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_17139_), .B(_17143_), .C(_17013_), .Y(_17144_) );
	NAND3X1 NAND3X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_17013_), .B(_17139_), .C(_17143_), .Y(_17145_) );
	INVX1 INVX1_1707 ( .gnd(gnd), .vdd(vdd), .A(_17145_), .Y(_17146_) );
	NOR2X1 NOR2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_17144_), .B(_17146_), .Y(_17147_) );
	OAI21X1 OAI21X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_16810_), .B(_17010_), .C(_17008_), .Y(_17148_) );
	XOR2X1 XOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_17147_), .B(_17148_), .Y(mulOut_11_) );
	AOI21X1 AOI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_17142_), .B(_17141_), .C(_17014_), .Y(_17149_) );
	AOI21X1 AOI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_17136_), .B(_17137_), .C(_16994_), .Y(_17150_) );
	INVX1 INVX1_1708 ( .gnd(gnd), .vdd(vdd), .A(_17129_), .Y(_17151_) );
	AOI21X1 AOI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_17118_), .B(_17112_), .C(_17021_), .Y(_17152_) );
	OAI21X1 OAI21X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_17018_), .B(_17152_), .C(_17119_), .Y(_17153_) );
	INVX1 INVX1_1709 ( .gnd(gnd), .vdd(vdd), .A(_17113_), .Y(_17154_) );
	AOI21X1 AOI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_17099_), .B(_17105_), .C(_17038_), .Y(_17155_) );
	OAI21X1 OAI21X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_17155_), .B(_17115_), .C(_17106_), .Y(_17156_) );
	INVX4 INVX4_14 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf2), .Y(_17157_) );
	NOR2X1 NOR2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf3), .B(_17157_), .Y(_17158_) );
	NAND2X1 NAND2X1_2495 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf1), .B(adder_bOperand_9_bF_buf3), .Y(_17159_) );
	NOR2X1 NOR2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_16876_), .B(_17159_), .Y(_17160_) );
	AOI21X1 AOI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_17026_), .B(_17023_), .C(_17160_), .Y(_17161_) );
	INVX1 INVX1_1710 ( .gnd(gnd), .vdd(vdd), .A(_17161_), .Y(_17162_) );
	NOR2X1 NOR2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_17022__bF_buf2), .Y(_17163_) );
	NAND2X1 NAND2X1_2496 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .B(adder_bOperand_9_bF_buf2), .Y(_17164_) );
	XOR2X1 XOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_17024_), .B(_17164_), .Y(_17165_) );
	NAND2X1 NAND2X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_17163_), .B(_17165_), .Y(_17166_) );
	NAND2X1 NAND2X1_2498 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(adder_bOperand_10_bF_buf1), .Y(_17167_) );
	OAI21X1 OAI21X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_17025__bF_buf2), .C(_17024_), .Y(_17168_) );
	OAI21X1 OAI21X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_17159_), .B(_17167_), .C(_17168_), .Y(_17169_) );
	OAI21X1 OAI21X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_17022__bF_buf1), .C(_17169_), .Y(_17170_) );
	NAND3X1 NAND3X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_17170_), .B(_17162_), .C(_17166_), .Y(_17171_) );
	INVX1 INVX1_1711 ( .gnd(gnd), .vdd(vdd), .A(_17163_), .Y(_17172_) );
	NOR2X1 NOR2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_17172_), .B(_17169_), .Y(_17173_) );
	INVX1 INVX1_1712 ( .gnd(gnd), .vdd(vdd), .A(_17170_), .Y(_17174_) );
	OAI21X1 OAI21X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_17173_), .B(_17174_), .C(_17161_), .Y(_17175_) );
	NAND3X1 NAND3X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_17158_), .B(_17171_), .C(_17175_), .Y(_17176_) );
	INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(_17158_), .Y(_17177_) );
	OAI21X1 OAI21X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_17173_), .B(_17174_), .C(_17162_), .Y(_17178_) );
	NAND3X1 NAND3X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_17161_), .B(_17170_), .C(_17166_), .Y(_17179_) );
	NAND3X1 NAND3X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_17177_), .B(_17179_), .C(_17178_), .Y(_17180_) );
	AOI21X1 AOI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_17046_), .B(_17047_), .C(_17051_), .Y(_17181_) );
	OAI21X1 OAI21X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_17041_), .B(_17181_), .C(_17052_), .Y(_17182_) );
	NAND3X1 NAND3X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_17182_), .B(_17176_), .C(_17180_), .Y(_17183_) );
	AOI21X1 AOI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_17178_), .B(_17179_), .C(_17177_), .Y(_17184_) );
	AOI21X1 AOI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_17175_), .B(_17171_), .C(_17158_), .Y(_17185_) );
	INVX1 INVX1_1713 ( .gnd(gnd), .vdd(vdd), .A(_17052_), .Y(_17186_) );
	AOI21X1 AOI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_17057_), .B(_17055_), .C(_17186_), .Y(_17187_) );
	OAI21X1 OAI21X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_17185_), .B(_17184_), .C(_17187_), .Y(_17188_) );
	NAND3X1 NAND3X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_17033_), .B(_17183_), .C(_17188_), .Y(_17189_) );
	NAND3X1 NAND3X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_17176_), .B(_17180_), .C(_17187_), .Y(_17190_) );
	OAI21X1 OAI21X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_17185_), .B(_17184_), .C(_17182_), .Y(_17191_) );
	NAND3X1 NAND3X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_17032_), .B(_17190_), .C(_17191_), .Y(_17192_) );
	NAND2X1 NAND2X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_17189_), .B(_17192_), .Y(_17193_) );
	AOI21X1 AOI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_17088_), .B(_17092_), .C(_17063_), .Y(_17194_) );
	OAI21X1 OAI21X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_17102_), .B(_17194_), .C(_17093_), .Y(_17195_) );
	OAI21X1 OAI21X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_17039_), .B(_17043_), .C(_17046_), .Y(_17196_) );
	NOR2X1 NOR2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf2), .B(_14728__bF_buf3), .Y(_17197_) );
	INVX1 INVX1_1714 ( .gnd(gnd), .vdd(vdd), .A(_17197_), .Y(_17198_) );
	NAND3X1 NAND3X1_2483 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf0), .B(adder_bOperand_6_bF_buf2), .C(_17043_), .Y(_17199_) );
	NAND2X1 NAND2X1_2500 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf4), .B(adder_bOperand_6_bF_buf1), .Y(_17200_) );
	NAND3X1 NAND3X1_2484 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf3), .B(adder_bOperand_7_bF_buf3), .C(_17200_), .Y(_17201_) );
	AOI21X1 AOI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_17199_), .B(_17201_), .C(_17198_), .Y(_17202_) );
	INVX1 INVX1_1715 ( .gnd(gnd), .vdd(vdd), .A(_17202_), .Y(_17203_) );
	NAND3X1 NAND3X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_17198_), .B(_17199_), .C(_17201_), .Y(_17204_) );
	NAND2X1 NAND2X1_2501 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf1), .B(aOperand_frameOut_8_bF_buf0), .Y(_17205_) );
	NOR2X1 NOR2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_16929_), .B(_17205_), .Y(_17206_) );
	AOI21X1 AOI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_17066_), .B(_17064_), .C(_17206_), .Y(_17207_) );
	INVX1 INVX1_1716 ( .gnd(gnd), .vdd(vdd), .A(_17207_), .Y(_17208_) );
	AOI21X1 AOI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_17203_), .B(_17204_), .C(_17208_), .Y(_17209_) );
	NAND2X1 NAND2X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_17199_), .B(_17201_), .Y(_17210_) );
	NOR2X1 NOR2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_17197_), .B(_17210_), .Y(_17211_) );
	NOR3X1 NOR3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_17207_), .B(_17202_), .C(_17211_), .Y(_17212_) );
	OAI21X1 OAI21X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_17212_), .B(_17209_), .C(_17196_), .Y(_17213_) );
	INVX1 INVX1_1717 ( .gnd(gnd), .vdd(vdd), .A(_17043_), .Y(_17214_) );
	AOI21X1 AOI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_17040_), .B(_17214_), .C(_17053_), .Y(_17215_) );
	OAI21X1 OAI21X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_17202_), .B(_17211_), .C(_17207_), .Y(_17216_) );
	NAND3X1 NAND3X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_17204_), .B(_17208_), .C(_17203_), .Y(_17217_) );
	NAND3X1 NAND3X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_17215_), .B(_17216_), .C(_17217_), .Y(_17218_) );
	NAND2X1 NAND2X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_17218_), .B(_17213_), .Y(_17219_) );
	AOI21X1 AOI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_17079_), .B(_17082_), .C(_17071_), .Y(_17220_) );
	OAI21X1 OAI21X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_17220_), .B(_17089_), .C(_17083_), .Y(_17221_) );
	NOR2X1 NOR2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf2), .B(_14049_), .Y(_17222_) );
	NAND2X1 NAND2X1_2504 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf1), .B(aOperand_frameOut_9_bF_buf0), .Y(_17223_) );
	OAI21X1 OAI21X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf0), .B(_15812__bF_buf3), .C(_17065_), .Y(_17224_) );
	OAI21X1 OAI21X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_17205_), .B(_17223_), .C(_17224_), .Y(_17225_) );
	OR2X2 OR2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_17225_), .B(_17222_), .Y(_17226_) );
	NAND2X1 NAND2X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_17222_), .B(_17225_), .Y(_17227_) );
	NAND2X1 NAND2X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_17227_), .B(_17226_), .Y(_17228_) );
	AOI21X1 AOI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_17078_), .B(_17073_), .C(_17080_), .Y(_17229_) );
	INVX1 INVX1_1718 ( .gnd(gnd), .vdd(vdd), .A(_17229_), .Y(_17230_) );
	NAND2X1 NAND2X1_2507 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf5), .B(aOperand_frameOut_10_bF_buf2), .Y(_17231_) );
	INVX1 INVX1_1719 ( .gnd(gnd), .vdd(vdd), .A(_17231_), .Y(_17232_) );
	NAND2X1 NAND2X1_2508 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf1), .B(aOperand_frameOut_11_bF_buf0), .Y(_17233_) );
	NAND2X1 NAND2X1_2509 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .B(aOperand_frameOut_12_bF_buf0), .Y(_17234_) );
	OR2X2 OR2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_17233_), .B(_17234_), .Y(_17235_) );
	INVX8 INVX8_68 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf4), .Y(_17236_) );
	OAI21X1 OAI21X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf2), .B(_17236__bF_buf3), .C(_17233_), .Y(_17237_) );
	NAND3X1 NAND3X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_17232_), .B(_17237_), .C(_17235_), .Y(_17238_) );
	NOR2X1 NOR2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_17233_), .B(_17234_), .Y(_17239_) );
	AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_17233_), .B(_17234_), .Y(_17240_) );
	OAI21X1 OAI21X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_17239_), .B(_17240_), .C(_17231_), .Y(_17241_) );
	NAND3X1 NAND3X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_17238_), .B(_17241_), .C(_17230_), .Y(_17242_) );
	NOR3X1 NOR3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_17231_), .B(_17239_), .C(_17240_), .Y(_17243_) );
	AOI21X1 AOI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_17235_), .B(_17237_), .C(_17232_), .Y(_17244_) );
	OAI21X1 OAI21X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_17244_), .B(_17243_), .C(_17229_), .Y(_17245_) );
	NAND3X1 NAND3X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_17245_), .B(_17242_), .C(_17228_), .Y(_17246_) );
	XOR2X1 XOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_17225_), .B(_17222_), .Y(_17247_) );
	OAI21X1 OAI21X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_17244_), .B(_17243_), .C(_17230_), .Y(_17248_) );
	NAND3X1 NAND3X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_17229_), .B(_17241_), .C(_17238_), .Y(_17249_) );
	NAND3X1 NAND3X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_17249_), .B(_17247_), .C(_17248_), .Y(_17250_) );
	NAND3X1 NAND3X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_17250_), .B(_17221_), .C(_17246_), .Y(_17251_) );
	INVX1 INVX1_1720 ( .gnd(gnd), .vdd(vdd), .A(_17083_), .Y(_17252_) );
	AOI21X1 AOI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_17087_), .B(_17070_), .C(_17252_), .Y(_17253_) );
	AOI21X1 AOI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_17248_), .B(_17249_), .C(_17247_), .Y(_17254_) );
	AOI21X1 AOI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_17242_), .B(_17245_), .C(_17228_), .Y(_17255_) );
	OAI21X1 OAI21X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_17254_), .B(_17255_), .C(_17253_), .Y(_17256_) );
	NAND3X1 NAND3X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_17251_), .B(_17256_), .C(_17219_), .Y(_17257_) );
	NAND3X1 NAND3X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_17216_), .B(_17196_), .C(_17217_), .Y(_17258_) );
	OAI21X1 OAI21X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_17212_), .B(_17209_), .C(_17215_), .Y(_17259_) );
	NAND2X1 NAND2X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_17258_), .B(_17259_), .Y(_17260_) );
	OAI21X1 OAI21X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_17254_), .B(_17255_), .C(_17221_), .Y(_17261_) );
	NAND3X1 NAND3X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_17250_), .B(_17246_), .C(_17253_), .Y(_17262_) );
	NAND3X1 NAND3X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_17262_), .B(_17261_), .C(_17260_), .Y(_17263_) );
	NAND3X1 NAND3X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_17195_), .B(_17257_), .C(_17263_), .Y(_17264_) );
	INVX1 INVX1_1721 ( .gnd(gnd), .vdd(vdd), .A(_17093_), .Y(_17265_) );
	AOI21X1 AOI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_17061_), .B(_17098_), .C(_17265_), .Y(_17266_) );
	AOI21X1 AOI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_17261_), .B(_17262_), .C(_17260_), .Y(_17267_) );
	AOI21X1 AOI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_17256_), .B(_17251_), .C(_17219_), .Y(_17268_) );
	OAI21X1 OAI21X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_17267_), .B(_17268_), .C(_17266_), .Y(_17269_) );
	NAND3X1 NAND3X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_17264_), .B(_17269_), .C(_17193_), .Y(_17270_) );
	NAND3X1 NAND3X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_17032_), .B(_17183_), .C(_17188_), .Y(_17271_) );
	NAND3X1 NAND3X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_17033_), .B(_17190_), .C(_17191_), .Y(_17272_) );
	NAND2X1 NAND2X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_17271_), .B(_17272_), .Y(_17273_) );
	OAI21X1 OAI21X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_17267_), .B(_17268_), .C(_17195_), .Y(_17274_) );
	NAND3X1 NAND3X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_17257_), .B(_17263_), .C(_17266_), .Y(_17275_) );
	NAND3X1 NAND3X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_17274_), .B(_17275_), .C(_17273_), .Y(_17276_) );
	NAND3X1 NAND3X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_17156_), .B(_17270_), .C(_17276_), .Y(_17277_) );
	INVX1 INVX1_1722 ( .gnd(gnd), .vdd(vdd), .A(_17106_), .Y(_17278_) );
	AOI21X1 AOI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_17036_), .B(_17111_), .C(_17278_), .Y(_17279_) );
	AOI22X1 AOI22X1_275 ( .gnd(gnd), .vdd(vdd), .A(_17189_), .B(_17192_), .C(_17274_), .D(_17275_), .Y(_17280_) );
	AOI21X1 AOI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_17269_), .B(_17264_), .C(_17193_), .Y(_17281_) );
	OAI21X1 OAI21X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_17280_), .B(_17281_), .C(_17279_), .Y(_17282_) );
	NAND3X1 NAND3X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_17154_), .B(_17277_), .C(_17282_), .Y(_17283_) );
	OAI21X1 OAI21X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_17280_), .B(_17281_), .C(_17156_), .Y(_17284_) );
	NAND3X1 NAND3X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_17270_), .B(_17276_), .C(_17279_), .Y(_17285_) );
	NAND3X1 NAND3X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_17113_), .B(_17285_), .C(_17284_), .Y(_17286_) );
	NAND3X1 NAND3X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_17153_), .B(_17283_), .C(_17286_), .Y(_17287_) );
	INVX1 INVX1_1723 ( .gnd(gnd), .vdd(vdd), .A(_17119_), .Y(_17288_) );
	AOI21X1 AOI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_17019_), .B(_17124_), .C(_17288_), .Y(_17289_) );
	AOI21X1 AOI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_17284_), .B(_17285_), .C(_17113_), .Y(_17290_) );
	AOI21X1 AOI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_17282_), .B(_17277_), .C(_17154_), .Y(_17291_) );
	OAI21X1 OAI21X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_17291_), .B(_17290_), .C(_17289_), .Y(_17292_) );
	NAND3X1 NAND3X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_17287_), .B(_17292_), .C(_17151_), .Y(_17293_) );
	OAI21X1 OAI21X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_17291_), .B(_17290_), .C(_17153_), .Y(_17294_) );
	NAND3X1 NAND3X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_17283_), .B(_17286_), .C(_17289_), .Y(_17296_) );
	NAND3X1 NAND3X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_17129_), .B(_17296_), .C(_17294_), .Y(_17297_) );
	NAND3X1 NAND3X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_17297_), .B(_17150_), .C(_17293_), .Y(_17298_) );
	AOI21X1 AOI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_17294_), .B(_17296_), .C(_17129_), .Y(_17299_) );
	NOR2X1 NOR2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_17133_), .B(_17132_), .Y(_17300_) );
	AOI22X1 AOI22X1_276 ( .gnd(gnd), .vdd(vdd), .A(_17017_), .B(_17300_), .C(_17287_), .D(_17292_), .Y(_17301_) );
	OAI21X1 OAI21X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_17301_), .B(_17299_), .C(_17135_), .Y(_17302_) );
	NAND3X1 NAND3X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_17149_), .B(_17298_), .C(_17302_), .Y(_17303_) );
	NAND3X1 NAND3X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_17140_), .B(_17135_), .C(_17138_), .Y(_17304_) );
	NAND3X1 NAND3X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_17135_), .B(_17297_), .C(_17293_), .Y(_17305_) );
	OAI21X1 OAI21X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_17301_), .B(_17299_), .C(_17150_), .Y(_17307_) );
	NAND3X1 NAND3X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_17304_), .B(_17305_), .C(_17307_), .Y(_17308_) );
	NAND2X1 NAND2X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_17303_), .B(_17308_), .Y(_17309_) );
	OAI21X1 OAI21X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_17144_), .B(_17148_), .C(_17145_), .Y(_17310_) );
	XOR2X1 XOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_17310_), .B(_17309_), .Y(mulOut_12_) );
	OAI21X1 OAI21X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_17309_), .B(_17310_), .C(_17303_), .Y(_17311_) );
	AOI21X1 AOI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_17276_), .B(_17270_), .C(_17156_), .Y(_17312_) );
	OAI21X1 OAI21X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_17113_), .B(_17312_), .C(_17277_), .Y(_17313_) );
	NAND2X1 NAND2X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_17183_), .B(_17271_), .Y(_17314_) );
	AOI21X1 AOI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_17257_), .B(_17263_), .C(_17195_), .Y(_17315_) );
	OAI21X1 OAI21X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_17315_), .B(_17273_), .C(_17264_), .Y(_17316_) );
	NAND2X1 NAND2X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_17171_), .B(_17176_), .Y(_17317_) );
	NAND2X1 NAND2X1_2515 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf2), .B(adder_bOperand_13_bF_buf0), .Y(_17318_) );
	INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf3), .Y(_17319_) );
	OAI22X1 OAI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf2), .B(_17319_), .C(_11874_), .D(_17157_), .Y(_17320_) );
	OAI21X1 OAI21X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_17318_), .B(_17177_), .C(_17320_), .Y(_17321_) );
	INVX1 INVX1_1724 ( .gnd(gnd), .vdd(vdd), .A(_17321_), .Y(_17322_) );
	NOR2X1 NOR2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_17024_), .B(_17164_), .Y(_17323_) );
	AOI21X1 AOI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_17168_), .B(_17163_), .C(_17323_), .Y(_17324_) );
	INVX1 INVX1_1725 ( .gnd(gnd), .vdd(vdd), .A(_17324_), .Y(_17325_) );
	NOR2X1 NOR2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf1), .B(_17022__bF_buf0), .Y(_11777_) );
	INVX1 INVX1_1726 ( .gnd(gnd), .vdd(vdd), .A(_11777_), .Y(_11778_) );
	NAND2X1 NAND2X1_2516 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .B(adder_bOperand_10_bF_buf0), .Y(_11779_) );
	OAI21X1 OAI21X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf1), .B(_17025__bF_buf1), .C(_17167_), .Y(_11780_) );
	OAI21X1 OAI21X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_17164_), .B(_11779_), .C(_11780_), .Y(_11781_) );
	OR2X2 OR2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_11781_), .B(_11778_), .Y(_11782_) );
	INVX1 INVX1_1727 ( .gnd(gnd), .vdd(vdd), .A(_17164_), .Y(_11783_) );
	INVX1 INVX1_1728 ( .gnd(gnd), .vdd(vdd), .A(_11779_), .Y(_11784_) );
	NAND2X1 NAND2X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_11783_), .B(_11784_), .Y(_11785_) );
	AOI21X1 AOI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_11785_), .B(_11780_), .C(_11777_), .Y(_11786_) );
	INVX1 INVX1_1729 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .Y(_11787_) );
	NAND3X1 NAND3X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_17325_), .B(_11782_), .C(_11787_), .Y(_11788_) );
	NOR2X1 NOR2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_11778_), .B(_11781_), .Y(_11789_) );
	OAI21X1 OAI21X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .B(_11789_), .C(_17324_), .Y(_11790_) );
	NAND3X1 NAND3X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_17322_), .B(_11790_), .C(_11788_), .Y(_11791_) );
	OAI21X1 OAI21X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .B(_11789_), .C(_17325_), .Y(_11792_) );
	NAND3X1 NAND3X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_17324_), .B(_11782_), .C(_11787_), .Y(_11793_) );
	NAND3X1 NAND3X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_17321_), .B(_11792_), .C(_11793_), .Y(_11794_) );
	OAI21X1 OAI21X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_17215_), .B(_17209_), .C(_17217_), .Y(_11795_) );
	NAND3X1 NAND3X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .B(_11794_), .C(_11795_), .Y(_11796_) );
	AOI21X1 AOI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_11793_), .B(_11792_), .C(_17321_), .Y(_11799_) );
	AOI21X1 AOI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_11788_), .B(_11790_), .C(_17322_), .Y(_11800_) );
	AOI21X1 AOI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_17196_), .B(_17216_), .C(_17212_), .Y(_11801_) );
	OAI21X1 OAI21X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_11799_), .B(_11800_), .C(_11801_), .Y(_11802_) );
	NAND3X1 NAND3X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_17317_), .B(_11796_), .C(_11802_), .Y(_11803_) );
	AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_17176_), .B(_17171_), .Y(_11804_) );
	NAND3X1 NAND3X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_11801_), .B(_11791_), .C(_11794_), .Y(_11805_) );
	OAI21X1 OAI21X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_11799_), .B(_11800_), .C(_11795_), .Y(_11806_) );
	NAND3X1 NAND3X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_11805_), .B(_11804_), .C(_11806_), .Y(_11807_) );
	AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_11807_), .B(_11803_), .Y(_11808_) );
	AOI21X1 AOI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_17246_), .B(_17250_), .C(_17221_), .Y(_11810_) );
	OAI21X1 OAI21X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_11810_), .B(_17260_), .C(_17251_), .Y(_11811_) );
	INVX1 INVX1_1730 ( .gnd(gnd), .vdd(vdd), .A(_17200_), .Y(_11812_) );
	AOI21X1 AOI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_17214_), .B(_11812_), .C(_17202_), .Y(_11813_) );
	INVX1 INVX1_1731 ( .gnd(gnd), .vdd(vdd), .A(_11813_), .Y(_11814_) );
	NOR2X1 NOR2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_14728__bF_buf2), .Y(_11815_) );
	INVX1 INVX1_1732 ( .gnd(gnd), .vdd(vdd), .A(_11815_), .Y(_11816_) );
	NAND2X1 NAND2X1_2518 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf3), .B(adder_bOperand_7_bF_buf2), .Y(_11817_) );
	NAND3X1 NAND3X1_2525 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf0), .B(aOperand_frameOut_7_bF_buf0), .C(_11817_), .Y(_11818_) );
	NAND2X1 NAND2X1_2519 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(aOperand_frameOut_7_bF_buf4), .Y(_11819_) );
	NAND3X1 NAND3X1_2526 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf2), .B(adder_bOperand_7_bF_buf1), .C(_11819_), .Y(_11821_) );
	AOI21X1 AOI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_11821_), .B(_11818_), .C(_11816_), .Y(_11822_) );
	NAND2X1 NAND2X1_2520 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf3), .B(adder_bOperand_7_bF_buf0), .Y(_11823_) );
	INVX1 INVX1_1733 ( .gnd(gnd), .vdd(vdd), .A(_11823_), .Y(_11824_) );
	NAND2X1 NAND2X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_11812_), .B(_11824_), .Y(_11825_) );
	OAI21X1 OAI21X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf3), .B(_14049_), .C(_11817_), .Y(_11826_) );
	AOI21X1 AOI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_11825_), .B(_11826_), .C(_11815_), .Y(_11827_) );
	NAND2X1 NAND2X1_2522 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf0), .B(aOperand_frameOut_9_bF_buf4), .Y(_11828_) );
	NOR2X1 NOR2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_17065_), .B(_11828_), .Y(_11829_) );
	AOI21X1 AOI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_17224_), .B(_17222_), .C(_11829_), .Y(_11830_) );
	OAI21X1 OAI21X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_11822_), .B(_11827_), .C(_11830_), .Y(_11832_) );
	NAND3X1 NAND3X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_11815_), .B(_11826_), .C(_11825_), .Y(_11833_) );
	NAND3X1 NAND3X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_11818_), .B(_11821_), .C(_11816_), .Y(_11834_) );
	INVX1 INVX1_1734 ( .gnd(gnd), .vdd(vdd), .A(_11830_), .Y(_11835_) );
	NAND3X1 NAND3X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11834_), .C(_11835_), .Y(_11836_) );
	NAND2X1 NAND2X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_11836_), .B(_11832_), .Y(_11837_) );
	XNOR2X1 XNOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_11837_), .B(_11814_), .Y(_11838_) );
	AOI21X1 AOI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_17238_), .B(_17241_), .C(_17230_), .Y(_11839_) );
	OAI21X1 OAI21X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_17247_), .B(_11839_), .C(_17242_), .Y(_11840_) );
	NOR2X1 NOR2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf1), .B(_15035_), .Y(_11841_) );
	NAND2X1 NAND2X1_2524 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf0), .B(aOperand_frameOut_10_bF_buf1), .Y(_11842_) );
	OAI21X1 OAI21X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf3), .B(_16940_), .C(_17223_), .Y(_11843_) );
	OAI21X1 OAI21X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_11828_), .B(_11842_), .C(_11843_), .Y(_11844_) );
	XNOR2X1 XNOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_11844_), .B(_11841_), .Y(_11845_) );
	AOI21X1 AOI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_17237_), .B(_17232_), .C(_17239_), .Y(_11846_) );
	INVX1 INVX1_1735 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .Y(_11847_) );
	NOR2X1 NOR2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_17077_), .Y(_11848_) );
	AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf0), .B(aOperand_frameOut_12_bF_buf3), .Y(_11849_) );
	AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(aOperand_frameOut_13_bF_buf0), .Y(_11850_) );
	NAND2X1 NAND2X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_11849_), .B(_11850_), .Y(_11851_) );
	NAND2X1 NAND2X1_2526 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .B(aOperand_frameOut_13_bF_buf4), .Y(_11853_) );
	OAI21X1 OAI21X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf1), .B(_17236__bF_buf2), .C(_11853_), .Y(_11854_) );
	NAND3X1 NAND3X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_11848_), .B(_11854_), .C(_11851_), .Y(_11855_) );
	INVX1 INVX1_1736 ( .gnd(gnd), .vdd(vdd), .A(_11848_), .Y(_11856_) );
	OAI21X1 OAI21X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf0), .B(_17236__bF_buf1), .C(_11850_), .Y(_11857_) );
	INVX4 INVX4_15 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf3), .Y(_11858_) );
	OAI21X1 OAI21X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf1), .B(_11858_), .C(_11849_), .Y(_11859_) );
	NAND3X1 NAND3X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_11857_), .B(_11859_), .C(_11856_), .Y(_11860_) );
	NAND3X1 NAND3X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_11855_), .B(_11860_), .C(_11847_), .Y(_11861_) );
	AOI21X1 AOI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_11857_), .B(_11859_), .C(_11856_), .Y(_11862_) );
	AOI21X1 AOI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_11851_), .B(_11854_), .C(_11848_), .Y(_11864_) );
	OAI21X1 OAI21X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_11864_), .B(_11862_), .C(_11846_), .Y(_11865_) );
	NAND3X1 NAND3X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_11845_), .B(_11865_), .C(_11861_), .Y(_11866_) );
	XOR2X1 XOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_11844_), .B(_11841_), .Y(_11867_) );
	OAI21X1 OAI21X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_11864_), .B(_11862_), .C(_11847_), .Y(_11868_) );
	NAND3X1 NAND3X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_11855_), .B(_11846_), .C(_11860_), .Y(_11869_) );
	NAND3X1 NAND3X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_11869_), .B(_11867_), .C(_11868_), .Y(_11870_) );
	NAND3X1 NAND3X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_11866_), .B(_11870_), .C(_11840_), .Y(_11871_) );
	INVX1 INVX1_1737 ( .gnd(gnd), .vdd(vdd), .A(_17242_), .Y(_11872_) );
	AOI21X1 AOI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_17228_), .B(_17245_), .C(_11872_), .Y(_11873_) );
	AOI21X1 AOI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_11868_), .B(_11869_), .C(_11867_), .Y(_11875_) );
	AOI21X1 AOI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_11861_), .B(_11865_), .C(_11845_), .Y(_11876_) );
	OAI21X1 OAI21X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_11875_), .B(_11876_), .C(_11873_), .Y(_11877_) );
	NAND3X1 NAND3X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_11871_), .B(_11877_), .C(_11838_), .Y(_11878_) );
	NAND3X1 NAND3X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_11832_), .B(_11836_), .C(_11814_), .Y(_11879_) );
	AOI21X1 AOI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11834_), .C(_11835_), .Y(_11880_) );
	NAND2X1 NAND2X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11834_), .Y(_11881_) );
	NOR2X1 NOR2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_11830_), .B(_11881_), .Y(_11882_) );
	OAI21X1 OAI21X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_11880_), .B(_11882_), .C(_11813_), .Y(_11883_) );
	NAND2X1 NAND2X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_11879_), .B(_11883_), .Y(_11884_) );
	OAI21X1 OAI21X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_11875_), .B(_11876_), .C(_11840_), .Y(_11886_) );
	NAND3X1 NAND3X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_11866_), .B(_11870_), .C(_11873_), .Y(_11887_) );
	NAND3X1 NAND3X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_11886_), .B(_11884_), .C(_11887_), .Y(_11888_) );
	NAND3X1 NAND3X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_11888_), .B(_11878_), .C(_11811_), .Y(_11889_) );
	INVX1 INVX1_1738 ( .gnd(gnd), .vdd(vdd), .A(_17251_), .Y(_11890_) );
	AOI21X1 AOI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_17219_), .B(_17256_), .C(_11890_), .Y(_11891_) );
	AOI21X1 AOI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_11886_), .C(_11884_), .Y(_11892_) );
	AOI21X1 AOI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_11877_), .B(_11871_), .C(_11838_), .Y(_11893_) );
	OAI21X1 OAI21X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_11893_), .B(_11892_), .C(_11891_), .Y(_11894_) );
	NAND3X1 NAND3X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_11889_), .B(_11894_), .C(_11808_), .Y(_11895_) );
	NAND2X1 NAND2X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_11803_), .B(_11807_), .Y(_11896_) );
	OAI21X1 OAI21X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_11893_), .B(_11892_), .C(_11811_), .Y(_11897_) );
	NAND3X1 NAND3X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_11888_), .B(_11878_), .C(_11891_), .Y(_11898_) );
	NAND3X1 NAND3X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_11896_), .B(_11898_), .C(_11897_), .Y(_11899_) );
	NAND3X1 NAND3X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_11899_), .B(_11895_), .C(_17316_), .Y(_11900_) );
	INVX1 INVX1_1739 ( .gnd(gnd), .vdd(vdd), .A(_17264_), .Y(_11901_) );
	AOI21X1 AOI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_17193_), .B(_17269_), .C(_11901_), .Y(_11902_) );
	AOI21X1 AOI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_11897_), .B(_11898_), .C(_11896_), .Y(_11903_) );
	AOI21X1 AOI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_11894_), .B(_11889_), .C(_11808_), .Y(_11904_) );
	OAI21X1 OAI21X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_11904_), .B(_11903_), .C(_11902_), .Y(_11905_) );
	NAND3X1 NAND3X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_17314_), .B(_11900_), .C(_11905_), .Y(_11907_) );
	INVX1 INVX1_1740 ( .gnd(gnd), .vdd(vdd), .A(_17314_), .Y(_11908_) );
	OAI21X1 OAI21X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_11904_), .B(_11903_), .C(_17316_), .Y(_11909_) );
	NAND3X1 NAND3X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_11895_), .B(_11899_), .C(_11902_), .Y(_11910_) );
	NAND3X1 NAND3X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_11908_), .B(_11910_), .C(_11909_), .Y(_11911_) );
	NAND3X1 NAND3X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_17313_), .B(_11907_), .C(_11911_), .Y(_11912_) );
	INVX1 INVX1_1741 ( .gnd(gnd), .vdd(vdd), .A(_17277_), .Y(_11913_) );
	AOI21X1 AOI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_17154_), .B(_17282_), .C(_11913_), .Y(_11914_) );
	AOI21X1 AOI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_11910_), .B(_11909_), .C(_11908_), .Y(_11915_) );
	AOI21X1 AOI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_11905_), .B(_11900_), .C(_17314_), .Y(_11916_) );
	OAI21X1 OAI21X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_11916_), .B(_11915_), .C(_11914_), .Y(_11919_) );
	NAND3X1 NAND3X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_17287_), .B(_11912_), .C(_11919_), .Y(_11920_) );
	INVX1 INVX1_1742 ( .gnd(gnd), .vdd(vdd), .A(_17287_), .Y(_11921_) );
	OAI21X1 OAI21X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_11916_), .B(_11915_), .C(_17313_), .Y(_11922_) );
	NAND3X1 NAND3X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_11907_), .B(_11911_), .C(_11914_), .Y(_11923_) );
	NAND3X1 NAND3X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_11923_), .B(_11922_), .C(_11921_), .Y(_11924_) );
	NAND2X1 NAND2X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_11920_), .B(_11924_), .Y(_11925_) );
	AOI21X1 AOI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_17150_), .B(_17297_), .C(_17299_), .Y(_11926_) );
	NAND2X1 NAND2X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_11925_), .B(_11926_), .Y(_11927_) );
	NAND3X1 NAND3X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_11912_), .B(_11919_), .C(_11921_), .Y(_11928_) );
	NAND3X1 NAND3X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_17287_), .B(_11923_), .C(_11922_), .Y(_11930_) );
	NAND2X1 NAND2X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_11930_), .B(_11928_), .Y(_11931_) );
	OAI21X1 OAI21X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_17135_), .B(_17301_), .C(_17293_), .Y(_11932_) );
	NAND2X1 NAND2X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_11931_), .B(_11932_), .Y(_11933_) );
	AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_11927_), .B(_11933_), .Y(_11934_) );
	XNOR2X1 XNOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_17311_), .B(_11934_), .Y(mulOut_13_) );
	INVX1 INVX1_1743 ( .gnd(gnd), .vdd(vdd), .A(_17298_), .Y(_11935_) );
	NAND2X1 NAND2X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_11925_), .B(_11935_), .Y(_11936_) );
	OAI21X1 OAI21X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_17303_), .B(_11934_), .C(_11936_), .Y(_11937_) );
	NOR3X1 NOR3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_11934_), .B(_17309_), .C(_17310_), .Y(_11938_) );
	NOR2X1 NOR2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_11937_), .B(_11938_), .Y(_11940_) );
	INVX1 INVX1_1744 ( .gnd(gnd), .vdd(vdd), .A(_11912_), .Y(_11941_) );
	AOI21X1 AOI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_11895_), .B(_11899_), .C(_17316_), .Y(_11942_) );
	OAI21X1 OAI21X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_11908_), .B(_11942_), .C(_11900_), .Y(_11943_) );
	OR2X2 OR2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_17177_), .B(_17318_), .Y(_11944_) );
	INVX1 INVX1_1745 ( .gnd(gnd), .vdd(vdd), .A(_11944_), .Y(_11945_) );
	NAND2X1 NAND2X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_11796_), .B(_11803_), .Y(_11946_) );
	XNOR2X1 XNOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_11946_), .B(_11945_), .Y(_11947_) );
	INVX1 INVX1_1746 ( .gnd(gnd), .vdd(vdd), .A(_11947_), .Y(_11948_) );
	AOI21X1 AOI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_11878_), .B(_11888_), .C(_11811_), .Y(_11949_) );
	OAI21X1 OAI21X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_11896_), .B(_11949_), .C(_11889_), .Y(_11951_) );
	AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .B(_11788_), .Y(_11952_) );
	NAND2X1 NAND2X1_2536 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf2), .B(adder_bOperand_14_bF_buf0), .Y(_11953_) );
	NAND2X1 NAND2X1_2537 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf0), .B(adder_bOperand_12_bF_buf1), .Y(_11954_) );
	XOR2X1 XOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_17318_), .B(_11954_), .Y(_11955_) );
	XNOR2X1 XNOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_11953_), .Y(_11956_) );
	AOI22X1 AOI22X1_277 ( .gnd(gnd), .vdd(vdd), .A(_11783_), .B(_11784_), .C(_11777_), .D(_11780_), .Y(_11957_) );
	INVX1 INVX1_1747 ( .gnd(gnd), .vdd(vdd), .A(_11957_), .Y(_11958_) );
	NOR2X1 NOR2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_17022__bF_buf3), .Y(_11959_) );
	INVX1 INVX1_1748 ( .gnd(gnd), .vdd(vdd), .A(_11959_), .Y(_11960_) );
	NAND2X1 NAND2X1_2538 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf2), .B(adder_bOperand_9_bF_buf1), .Y(_11961_) );
	NAND2X1 NAND2X1_2539 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf2), .B(adder_bOperand_10_bF_buf4), .Y(_11962_) );
	OAI21X1 OAI21X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_17025__bF_buf0), .C(_11779_), .Y(_11963_) );
	OAI21X1 OAI21X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_11961_), .B(_11962_), .C(_11963_), .Y(_11964_) );
	OR2X2 OR2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_11964_), .B(_11960_), .Y(_11965_) );
	OAI21X1 OAI21X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_17022__bF_buf2), .C(_11964_), .Y(_11966_) );
	NAND3X1 NAND3X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_11966_), .B(_11958_), .C(_11965_), .Y(_11967_) );
	NOR2X1 NOR2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_11960_), .B(_11964_), .Y(_11968_) );
	NAND2X1 NAND2X1_2540 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf1), .B(adder_bOperand_9_bF_buf0), .Y(_11969_) );
	NOR2X1 NOR2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_11779_), .B(_11969_), .Y(_11970_) );
	INVX1 INVX1_1749 ( .gnd(gnd), .vdd(vdd), .A(_11970_), .Y(_11972_) );
	AOI21X1 AOI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_11972_), .B(_11963_), .C(_11959_), .Y(_11973_) );
	OAI21X1 OAI21X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_11968_), .B(_11973_), .C(_11957_), .Y(_11974_) );
	NAND3X1 NAND3X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_11956_), .B(_11974_), .C(_11967_), .Y(_11975_) );
	XOR2X1 XOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_11953_), .Y(_11976_) );
	OAI21X1 OAI21X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_11968_), .B(_11973_), .C(_11958_), .Y(_11977_) );
	NAND3X1 NAND3X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_11957_), .B(_11966_), .C(_11965_), .Y(_11978_) );
	NAND3X1 NAND3X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_11976_), .B(_11977_), .C(_11978_), .Y(_11979_) );
	OAI21X1 OAI21X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_11813_), .B(_11880_), .C(_11836_), .Y(_11980_) );
	NAND3X1 NAND3X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_11980_), .B(_11975_), .C(_11979_), .Y(_11981_) );
	AOI21X1 AOI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_11978_), .B(_11977_), .C(_11976_), .Y(_11983_) );
	AOI21X1 AOI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_11967_), .B(_11974_), .C(_11956_), .Y(_11984_) );
	INVX1 INVX1_1750 ( .gnd(gnd), .vdd(vdd), .A(_11980_), .Y(_11985_) );
	OAI21X1 OAI21X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_11984_), .C(_11985_), .Y(_11986_) );
	NAND3X1 NAND3X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_11981_), .B(_11952_), .C(_11986_), .Y(_11987_) );
	NAND2X1 NAND2X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_11788_), .B(_11791_), .Y(_11988_) );
	NAND3X1 NAND3X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_11975_), .B(_11979_), .C(_11985_), .Y(_11989_) );
	OAI21X1 OAI21X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_11984_), .C(_11980_), .Y(_11990_) );
	NAND3X1 NAND3X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_11988_), .B(_11990_), .C(_11989_), .Y(_11991_) );
	NAND2X1 NAND2X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_11987_), .B(_11991_), .Y(_11992_) );
	AOI21X1 AOI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_11866_), .B(_11870_), .C(_11840_), .Y(_11994_) );
	OAI21X1 OAI21X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_11994_), .B(_11884_), .C(_11871_), .Y(_11995_) );
	OAI21X1 OAI21X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_17200_), .B(_11823_), .C(_11833_), .Y(_11996_) );
	INVX1 INVX1_1751 ( .gnd(gnd), .vdd(vdd), .A(_11996_), .Y(_11997_) );
	NOR2X1 NOR2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf0), .B(_14728__bF_buf1), .Y(_11998_) );
	NAND2X1 NAND2X1_2543 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf4), .B(aOperand_frameOut_8_bF_buf4), .Y(_11999_) );
	INVX1 INVX1_1752 ( .gnd(gnd), .vdd(vdd), .A(_11999_), .Y(_12000_) );
	NAND2X1 NAND2X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_11824_), .B(_12000_), .Y(_12001_) );
	OAI21X1 OAI21X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf2), .B(_15035_), .C(_11823_), .Y(_12002_) );
	NAND3X1 NAND3X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_11998_), .B(_12002_), .C(_12001_), .Y(_12003_) );
	NAND2X1 NAND2X1_2545 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(aOperand_frameOut_8_bF_buf3), .Y(_12005_) );
	OAI21X1 OAI21X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_11819_), .B(_12005_), .C(_12002_), .Y(_12006_) );
	OAI21X1 OAI21X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf3), .B(_14728__bF_buf0), .C(_12006_), .Y(_12007_) );
	NAND2X1 NAND2X1_2546 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf5), .B(aOperand_frameOut_10_bF_buf0), .Y(_12008_) );
	NOR2X1 NOR2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_17223_), .B(_12008_), .Y(_12009_) );
	AOI21X1 AOI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_11843_), .B(_11841_), .C(_12009_), .Y(_12010_) );
	INVX1 INVX1_1753 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .Y(_12011_) );
	NAND3X1 NAND3X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_12003_), .B(_12007_), .C(_12011_), .Y(_12012_) );
	INVX1 INVX1_1754 ( .gnd(gnd), .vdd(vdd), .A(_12003_), .Y(_12013_) );
	AOI21X1 AOI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .B(_12002_), .C(_11998_), .Y(_12014_) );
	OAI21X1 OAI21X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_12014_), .B(_12013_), .C(_12010_), .Y(_12016_) );
	NAND3X1 NAND3X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_11997_), .B(_12012_), .C(_12016_), .Y(_12017_) );
	NAND3X1 NAND3X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .B(_12003_), .C(_12007_), .Y(_12018_) );
	OAI21X1 OAI21X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_12014_), .B(_12013_), .C(_12011_), .Y(_12019_) );
	NAND3X1 NAND3X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_11996_), .B(_12018_), .C(_12019_), .Y(_12020_) );
	NAND2X1 NAND2X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_12020_), .B(_12017_), .Y(_12021_) );
	AOI21X1 AOI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .B(_11855_), .C(_11847_), .Y(_12022_) );
	OAI21X1 OAI21X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_11867_), .B(_12022_), .C(_11861_), .Y(_12023_) );
	NOR2X1 NOR2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf0), .B(_15812__bF_buf2), .Y(_12024_) );
	NAND2X1 NAND2X1_2548 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf5), .B(aOperand_frameOut_11_bF_buf4), .Y(_12025_) );
	OAI21X1 OAI21X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf2), .B(_17077_), .C(_11842_), .Y(_12027_) );
	OAI21X1 OAI21X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_12008_), .B(_12025_), .C(_12027_), .Y(_12028_) );
	XNOR2X1 XNOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_12028_), .B(_12024_), .Y(_12029_) );
	INVX1 INVX1_1755 ( .gnd(gnd), .vdd(vdd), .A(_17234_), .Y(_12030_) );
	AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf6), .B(aOperand_frameOut_13_bF_buf2), .Y(_12031_) );
	AOI22X1 AOI22X1_278 ( .gnd(gnd), .vdd(vdd), .A(_12030_), .B(_12031_), .C(_11848_), .D(_11854_), .Y(_12032_) );
	INVX1 INVX1_1756 ( .gnd(gnd), .vdd(vdd), .A(_12032_), .Y(_12033_) );
	NAND2X1 NAND2X1_2549 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .B(aOperand_frameOut_12_bF_buf2), .Y(_12034_) );
	INVX1 INVX1_1757 ( .gnd(gnd), .vdd(vdd), .A(_12034_), .Y(_12035_) );
	AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_14_bF_buf1), .Y(_12036_) );
	NAND2X1 NAND2X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_12031_), .B(_12036_), .Y(_12038_) );
	INVX4 INVX4_16 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf0), .Y(_12039_) );
	OAI22X1 OAI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf0), .B(_12039_), .C(_11776__bF_buf3), .D(_11858_), .Y(_12040_) );
	NAND3X1 NAND3X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_12035_), .B(_12040_), .C(_12038_), .Y(_12041_) );
	NAND2X1 NAND2X1_2551 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(aOperand_frameOut_14_bF_buf4), .Y(_12042_) );
	NOR2X1 NOR2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_11853_), .B(_12042_), .Y(_12043_) );
	NOR2X1 NOR2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_12031_), .B(_12036_), .Y(_12044_) );
	OAI21X1 OAI21X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_12043_), .B(_12044_), .C(_12034_), .Y(_12045_) );
	NAND3X1 NAND3X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_12041_), .B(_12045_), .C(_12033_), .Y(_12046_) );
	OAI21X1 OAI21X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf2), .B(_11858_), .C(_12036_), .Y(_12047_) );
	OAI21X1 OAI21X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf4), .B(_12039_), .C(_12031_), .Y(_12049_) );
	AOI21X1 AOI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_12047_), .B(_12049_), .C(_12034_), .Y(_12050_) );
	AOI21X1 AOI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_12038_), .B(_12040_), .C(_12035_), .Y(_12051_) );
	OAI21X1 OAI21X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_12051_), .B(_12050_), .C(_12032_), .Y(_12052_) );
	NAND3X1 NAND3X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_12052_), .B(_12029_), .C(_12046_), .Y(_12053_) );
	XOR2X1 XOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_12028_), .B(_12024_), .Y(_12054_) );
	NOR3X1 NOR3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_12032_), .B(_12051_), .C(_12050_), .Y(_12055_) );
	AOI21X1 AOI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_12045_), .B(_12041_), .C(_12033_), .Y(_12056_) );
	OAI21X1 OAI21X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_12056_), .B(_12055_), .C(_12054_), .Y(_12057_) );
	NAND3X1 NAND3X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_12053_), .B(_12023_), .C(_12057_), .Y(_12058_) );
	NOR3X1 NOR3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .B(_11864_), .C(_11862_), .Y(_12060_) );
	AOI21X1 AOI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_11865_), .B(_11845_), .C(_12060_), .Y(_12061_) );
	OAI21X1 OAI21X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_12051_), .B(_12050_), .C(_12033_), .Y(_12062_) );
	NAND3X1 NAND3X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_12032_), .B(_12041_), .C(_12045_), .Y(_12063_) );
	AOI21X1 AOI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_12062_), .B(_12063_), .C(_12054_), .Y(_12064_) );
	AOI21X1 AOI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_12046_), .B(_12052_), .C(_12029_), .Y(_12065_) );
	OAI21X1 OAI21X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_12064_), .B(_12065_), .C(_12061_), .Y(_12066_) );
	NAND3X1 NAND3X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_12058_), .B(_12021_), .C(_12066_), .Y(_12067_) );
	NAND3X1 NAND3X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_11996_), .B(_12012_), .C(_12016_), .Y(_12068_) );
	NAND3X1 NAND3X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_11997_), .B(_12018_), .C(_12019_), .Y(_12069_) );
	NAND2X1 NAND2X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_12069_), .B(_12068_), .Y(_12071_) );
	OAI21X1 OAI21X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_12064_), .B(_12065_), .C(_12023_), .Y(_12072_) );
	NAND3X1 NAND3X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_12053_), .B(_12061_), .C(_12057_), .Y(_12073_) );
	NAND3X1 NAND3X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_12073_), .B(_12072_), .C(_12071_), .Y(_12074_) );
	NAND3X1 NAND3X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_12067_), .B(_12074_), .C(_11995_), .Y(_12075_) );
	INVX1 INVX1_1758 ( .gnd(gnd), .vdd(vdd), .A(_11871_), .Y(_12076_) );
	AOI21X1 AOI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_11838_), .B(_11877_), .C(_12076_), .Y(_12077_) );
	AOI21X1 AOI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_12072_), .B(_12073_), .C(_12071_), .Y(_12078_) );
	AOI21X1 AOI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_12066_), .B(_12058_), .C(_12021_), .Y(_12079_) );
	OAI21X1 OAI21X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_12078_), .B(_12079_), .C(_12077_), .Y(_12080_) );
	NAND3X1 NAND3X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_12075_), .B(_11992_), .C(_12080_), .Y(_12082_) );
	NAND3X1 NAND3X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_11988_), .B(_11981_), .C(_11986_), .Y(_12083_) );
	NAND3X1 NAND3X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_11952_), .B(_11990_), .C(_11989_), .Y(_12084_) );
	NAND2X1 NAND2X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_12083_), .B(_12084_), .Y(_12085_) );
	OAI21X1 OAI21X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_12078_), .B(_12079_), .C(_11995_), .Y(_12086_) );
	NAND3X1 NAND3X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_12067_), .B(_12074_), .C(_12077_), .Y(_12087_) );
	NAND3X1 NAND3X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_12085_), .B(_12086_), .C(_12087_), .Y(_12088_) );
	NAND3X1 NAND3X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_12088_), .C(_11951_), .Y(_12089_) );
	INVX1 INVX1_1759 ( .gnd(gnd), .vdd(vdd), .A(_11889_), .Y(_12090_) );
	AOI21X1 AOI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_11808_), .B(_11894_), .C(_12090_), .Y(_12091_) );
	AOI21X1 AOI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_12087_), .B(_12086_), .C(_12085_), .Y(_12093_) );
	AOI21X1 AOI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_12080_), .B(_12075_), .C(_11992_), .Y(_12094_) );
	OAI21X1 OAI21X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_12094_), .B(_12093_), .C(_12091_), .Y(_12095_) );
	NAND3X1 NAND3X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_12089_), .B(_11948_), .C(_12095_), .Y(_12096_) );
	INVX1 INVX1_1760 ( .gnd(gnd), .vdd(vdd), .A(_12089_), .Y(_12097_) );
	AOI21X1 AOI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_12088_), .B(_12082_), .C(_11951_), .Y(_12098_) );
	OAI21X1 OAI21X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_12098_), .B(_12097_), .C(_11947_), .Y(_12099_) );
	NAND3X1 NAND3X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_11943_), .B(_12096_), .C(_12099_), .Y(_12100_) );
	INVX1 INVX1_1761 ( .gnd(gnd), .vdd(vdd), .A(_11900_), .Y(_12101_) );
	AOI21X1 AOI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_17314_), .B(_11905_), .C(_12101_), .Y(_12102_) );
	OAI21X1 OAI21X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_12094_), .B(_12093_), .C(_11951_), .Y(_12104_) );
	NAND3X1 NAND3X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_12088_), .C(_12091_), .Y(_12105_) );
	AOI21X1 AOI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_12105_), .B(_12104_), .C(_11947_), .Y(_12106_) );
	AOI21X1 AOI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_12095_), .B(_12089_), .C(_11948_), .Y(_12107_) );
	OAI21X1 OAI21X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_12107_), .B(_12106_), .C(_12102_), .Y(_12108_) );
	NAND3X1 NAND3X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_12100_), .B(_12108_), .C(_11941_), .Y(_12109_) );
	OAI21X1 OAI21X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_12107_), .B(_12106_), .C(_11943_), .Y(_12110_) );
	NAND3X1 NAND3X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_12096_), .B(_12099_), .C(_12102_), .Y(_12111_) );
	NAND3X1 NAND3X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_11912_), .B(_12110_), .C(_12111_), .Y(_12112_) );
	NAND2X1 NAND2X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_12112_), .B(_12109_), .Y(_12113_) );
	AOI21X1 AOI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_11919_), .B(_11912_), .C(_11921_), .Y(_12115_) );
	OAI21X1 OAI21X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_17293_), .B(_12115_), .C(_11928_), .Y(_12116_) );
	NOR2X1 NOR2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_12113_), .B(_12116_), .Y(_12117_) );
	INVX1 INVX1_1762 ( .gnd(gnd), .vdd(vdd), .A(_12117_), .Y(_12118_) );
	AOI21X1 AOI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_12111_), .B(_12110_), .C(_11912_), .Y(_12119_) );
	NOR2X1 NOR2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_11916_), .B(_11915_), .Y(_12120_) );
	AOI22X1 AOI22X1_279 ( .gnd(gnd), .vdd(vdd), .A(_12120_), .B(_17313_), .C(_12108_), .D(_12100_), .Y(_12121_) );
	OAI21X1 OAI21X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_12119_), .B(_12121_), .C(_12116_), .Y(_12122_) );
	NAND2X1 NAND2X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_12122_), .B(_12118_), .Y(_12123_) );
	XNOR2X1 XNOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_11940_), .B(_12123_), .Y(mulOut_14_) );
	NAND3X1 NAND3X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_17299_), .B(_11930_), .C(_11928_), .Y(_12125_) );
	OAI21X1 OAI21X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_11937_), .B(_11938_), .C(_12123_), .Y(_12126_) );
	OAI21X1 OAI21X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_12113_), .B(_12125_), .C(_12126_), .Y(_12127_) );
	INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(_12100_), .Y(_12128_) );
	NAND2X1 NAND2X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_11945_), .B(_11946_), .Y(_12129_) );
	OAI21X1 OAI21X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_11947_), .B(_12098_), .C(_12089_), .Y(_12130_) );
	INVX8 INVX8_69 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf0), .Y(_12131_) );
	NOR2X1 NOR2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf1), .B(_12131_), .Y(_12132_) );
	NAND3X1 NAND3X1_2592 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf1), .B(adder_bOperand_14_bF_buf3), .C(_11955_), .Y(_12133_) );
	OAI21X1 OAI21X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_17318_), .B(_11954_), .C(_12133_), .Y(_12134_) );
	NOR2X1 NOR2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .B(_12134_), .Y(_12136_) );
	NAND2X1 NAND2X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_12132_), .B(_12134_), .Y(_12137_) );
	INVX1 INVX1_1763 ( .gnd(gnd), .vdd(vdd), .A(_12137_), .Y(_12138_) );
	NOR2X1 NOR2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_12136_), .B(_12138_), .Y(_12139_) );
	NAND2X1 NAND2X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_11981_), .B(_12083_), .Y(_12140_) );
	NAND2X1 NAND2X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_12139_), .B(_12140_), .Y(_12141_) );
	OR2X2 OR2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_12140_), .B(_12139_), .Y(_12142_) );
	AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_12142_), .B(_12141_), .Y(_12143_) );
	AOI21X1 AOI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_12067_), .B(_12074_), .C(_11995_), .Y(_12144_) );
	OAI21X1 OAI21X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_12085_), .B(_12144_), .C(_12075_), .Y(_12145_) );
	AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_11975_), .B(_11967_), .Y(_12147_) );
	NAND2X1 NAND2X1_2560 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf1), .B(adder_bOperand_14_bF_buf2), .Y(_12148_) );
	NAND2X1 NAND2X1_2561 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf0), .B(adder_bOperand_13_bF_buf2), .Y(_12149_) );
	NAND2X1 NAND2X1_2562 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf4), .B(adder_bOperand_12_bF_buf0), .Y(_12150_) );
	OAI21X1 OAI21X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf0), .B(_17319_), .C(_12150_), .Y(_12151_) );
	OAI21X1 OAI21X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_12149_), .C(_12151_), .Y(_12152_) );
	XOR2X1 XOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_12152_), .B(_12148_), .Y(_12153_) );
	AOI21X1 AOI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_11963_), .B(_11959_), .C(_11970_), .Y(_12154_) );
	INVX1 INVX1_1764 ( .gnd(gnd), .vdd(vdd), .A(_12154_), .Y(_12155_) );
	NOR2X1 NOR2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf0), .B(_17022__bF_buf1), .Y(_12156_) );
	INVX1 INVX1_1765 ( .gnd(gnd), .vdd(vdd), .A(_12156_), .Y(_12158_) );
	NAND2X1 NAND2X1_2563 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf1), .B(adder_bOperand_10_bF_buf3), .Y(_12159_) );
	OAI21X1 OAI21X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf2), .B(_17025__bF_buf3), .C(_11962_), .Y(_12160_) );
	OAI21X1 OAI21X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_11969_), .B(_12159_), .C(_12160_), .Y(_12161_) );
	OR2X2 OR2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_12161_), .B(_12158_), .Y(_12162_) );
	OAI21X1 OAI21X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf3), .B(_17022__bF_buf0), .C(_12161_), .Y(_12163_) );
	NAND3X1 NAND3X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_12163_), .B(_12155_), .C(_12162_), .Y(_12164_) );
	NOR2X1 NOR2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_12158_), .B(_12161_), .Y(_12165_) );
	INVX1 INVX1_1766 ( .gnd(gnd), .vdd(vdd), .A(_11969_), .Y(_12166_) );
	INVX1 INVX1_1767 ( .gnd(gnd), .vdd(vdd), .A(_12159_), .Y(_12167_) );
	NAND2X1 NAND2X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_12166_), .B(_12167_), .Y(_12168_) );
	AOI21X1 AOI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_12168_), .B(_12160_), .C(_12156_), .Y(_12169_) );
	OAI21X1 OAI21X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_12169_), .B(_12165_), .C(_12154_), .Y(_12170_) );
	NAND3X1 NAND3X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_12153_), .B(_12170_), .C(_12164_), .Y(_12171_) );
	INVX1 INVX1_1768 ( .gnd(gnd), .vdd(vdd), .A(_12153_), .Y(_12172_) );
	OAI21X1 OAI21X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_12169_), .B(_12165_), .C(_12155_), .Y(_12173_) );
	NAND3X1 NAND3X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_12154_), .B(_12163_), .C(_12162_), .Y(_12174_) );
	NAND3X1 NAND3X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_12173_), .B(_12174_), .C(_12172_), .Y(_12175_) );
	AOI21X1 AOI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_12007_), .B(_12003_), .C(_12011_), .Y(_12176_) );
	OAI21X1 OAI21X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_12176_), .B(_11997_), .C(_12012_), .Y(_12177_) );
	NAND3X1 NAND3X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_12171_), .B(_12177_), .C(_12175_), .Y(_12180_) );
	AOI21X1 AOI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_12174_), .B(_12173_), .C(_12172_), .Y(_12181_) );
	AOI21X1 AOI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_12164_), .B(_12170_), .C(_12153_), .Y(_12182_) );
	INVX1 INVX1_1769 ( .gnd(gnd), .vdd(vdd), .A(_12177_), .Y(_12183_) );
	OAI21X1 OAI21X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_12181_), .B(_12182_), .C(_12183_), .Y(_12184_) );
	NAND3X1 NAND3X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_12147_), .B(_12180_), .C(_12184_), .Y(_12185_) );
	NAND2X1 NAND2X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_11967_), .B(_11975_), .Y(_12186_) );
	NAND3X1 NAND3X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_12171_), .B(_12175_), .C(_12183_), .Y(_12187_) );
	OAI21X1 OAI21X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_12182_), .B(_12181_), .C(_12177_), .Y(_12188_) );
	NAND3X1 NAND3X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_12186_), .B(_12188_), .C(_12187_), .Y(_12189_) );
	NAND2X1 NAND2X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_12185_), .B(_12189_), .Y(_12191_) );
	AOI21X1 AOI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_12057_), .B(_12053_), .C(_12023_), .Y(_12192_) );
	OAI21X1 OAI21X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_12071_), .B(_12192_), .C(_12058_), .Y(_12193_) );
	OAI21X1 OAI21X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_11819_), .B(_12005_), .C(_12003_), .Y(_12194_) );
	NAND2X1 NAND2X1_2567 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf2), .B(adder_bOperand_8_bF_buf0), .Y(_12195_) );
	NAND2X1 NAND2X1_2568 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf4), .B(aOperand_frameOut_9_bF_buf3), .Y(_12196_) );
	OAI21X1 OAI21X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf1), .B(_15812__bF_buf1), .C(_12005_), .Y(_12197_) );
	OAI21X1 OAI21X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_11999_), .B(_12196_), .C(_12197_), .Y(_12198_) );
	OR2X2 OR2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_12198_), .B(_12195_), .Y(_12199_) );
	OAI21X1 OAI21X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_14728__bF_buf3), .C(_12198_), .Y(_12200_) );
	NAND2X1 NAND2X1_2569 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .B(aOperand_frameOut_11_bF_buf3), .Y(_12202_) );
	NOR2X1 NOR2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_11842_), .B(_12202_), .Y(_12203_) );
	AOI21X1 AOI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_12027_), .B(_12024_), .C(_12203_), .Y(_12204_) );
	INVX1 INVX1_1770 ( .gnd(gnd), .vdd(vdd), .A(_12204_), .Y(_12205_) );
	NAND3X1 NAND3X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12205_), .C(_12199_), .Y(_12206_) );
	NOR2X1 NOR2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_12195_), .B(_12198_), .Y(_12207_) );
	INVX1 INVX1_1771 ( .gnd(gnd), .vdd(vdd), .A(_12196_), .Y(_12208_) );
	NAND2X1 NAND2X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_12000_), .B(_12208_), .Y(_12209_) );
	AOI22X1 AOI22X1_280 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf1), .B(adder_bOperand_8_bF_buf4), .C(_12197_), .D(_12209_), .Y(_12210_) );
	OAI21X1 OAI21X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_12210_), .B(_12207_), .C(_12204_), .Y(_12211_) );
	NAND3X1 NAND3X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_12194_), .B(_12211_), .C(_12206_), .Y(_12213_) );
	INVX1 INVX1_1772 ( .gnd(gnd), .vdd(vdd), .A(_12194_), .Y(_12214_) );
	NAND3X1 NAND3X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12204_), .C(_12199_), .Y(_12215_) );
	OAI21X1 OAI21X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_12210_), .B(_12207_), .C(_12205_), .Y(_12216_) );
	NAND3X1 NAND3X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_12216_), .B(_12214_), .C(_12215_), .Y(_12217_) );
	AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_12217_), .B(_12213_), .Y(_12218_) );
	OAI21X1 OAI21X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_12054_), .B(_12056_), .C(_12046_), .Y(_12219_) );
	NAND2X1 NAND2X1_2571 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf0), .B(aOperand_frameOut_10_bF_buf4), .Y(_12220_) );
	INVX1 INVX1_1773 ( .gnd(gnd), .vdd(vdd), .A(_12220_), .Y(_12221_) );
	NAND2X1 NAND2X1_2572 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .B(aOperand_frameOut_12_bF_buf1), .Y(_12222_) );
	OAI21X1 OAI21X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf1), .B(_17236__bF_buf0), .C(_12025_), .Y(_12224_) );
	OAI21X1 OAI21X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_12202_), .B(_12222_), .C(_12224_), .Y(_12225_) );
	XNOR2X1 XNOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_12225_), .B(_12221_), .Y(_12226_) );
	OAI21X1 OAI21X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_12034_), .B(_12044_), .C(_12038_), .Y(_12227_) );
	NAND2X1 NAND2X1_2573 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf3), .B(aOperand_frameOut_13_bF_buf1), .Y(_12228_) );
	INVX1 INVX1_1774 ( .gnd(gnd), .vdd(vdd), .A(_12228_), .Y(_12229_) );
	AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf4), .B(aOperand_frameOut_14_bF_buf3), .Y(_12230_) );
	AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_15_bF_buf1), .Y(_12231_) );
	NAND2X1 NAND2X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_12230_), .B(_12231_), .Y(_12232_) );
	INVX8 INVX8_70 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf0), .Y(_12233_) );
	OAI21X1 OAI21X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf3), .B(_12233_), .C(_12042_), .Y(_12234_) );
	NAND3X1 NAND3X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_12229_), .B(_12234_), .C(_12232_), .Y(_12235_) );
	NAND2X1 NAND2X1_2575 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_15_bF_buf4), .Y(_12236_) );
	NOR2X1 NOR2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_12042_), .B(_12236_), .Y(_12237_) );
	AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_12042_), .B(_12236_), .Y(_12238_) );
	OAI21X1 OAI21X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_12237_), .B(_12238_), .C(_12228_), .Y(_12239_) );
	NAND3X1 NAND3X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_12235_), .B(_12239_), .C(_12227_), .Y(_12240_) );
	AOI21X1 AOI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_12040_), .B(_12035_), .C(_12043_), .Y(_12241_) );
	OAI21X1 OAI21X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf1), .B(_12039_), .C(_12231_), .Y(_12242_) );
	OAI21X1 OAI21X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf2), .B(_12233_), .C(_12230_), .Y(_12243_) );
	AOI21X1 AOI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_12242_), .B(_12243_), .C(_12228_), .Y(_12245_) );
	AOI21X1 AOI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_12232_), .B(_12234_), .C(_12229_), .Y(_12246_) );
	OAI21X1 OAI21X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_12246_), .B(_12245_), .C(_12241_), .Y(_12247_) );
	NAND3X1 NAND3X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_12240_), .B(_12247_), .C(_12226_), .Y(_12248_) );
	XNOR2X1 XNOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_12225_), .B(_12220_), .Y(_12249_) );
	OAI21X1 OAI21X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_12246_), .B(_12245_), .C(_12227_), .Y(_12250_) );
	NAND3X1 NAND3X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_12235_), .B(_12241_), .C(_12239_), .Y(_12251_) );
	NAND3X1 NAND3X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_12251_), .B(_12250_), .C(_12249_), .Y(_12252_) );
	NAND3X1 NAND3X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_12248_), .B(_12252_), .C(_12219_), .Y(_12253_) );
	AOI21X1 AOI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_12029_), .B(_12052_), .C(_12055_), .Y(_12254_) );
	AOI21X1 AOI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_12250_), .B(_12251_), .C(_12249_), .Y(_12256_) );
	AOI21X1 AOI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_12247_), .B(_12240_), .C(_12226_), .Y(_12257_) );
	OAI21X1 OAI21X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_12256_), .B(_12257_), .C(_12254_), .Y(_12258_) );
	NAND3X1 NAND3X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_12253_), .B(_12258_), .C(_12218_), .Y(_12259_) );
	NAND2X1 NAND2X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_12213_), .B(_12217_), .Y(_12260_) );
	OAI21X1 OAI21X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_12256_), .B(_12257_), .C(_12219_), .Y(_12261_) );
	NAND3X1 NAND3X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_12248_), .B(_12252_), .C(_12254_), .Y(_12262_) );
	NAND3X1 NAND3X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_12262_), .B(_12261_), .C(_12260_), .Y(_12263_) );
	NAND3X1 NAND3X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_12263_), .B(_12259_), .C(_12193_), .Y(_12264_) );
	NOR3X1 NOR3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_12064_), .B(_12065_), .C(_12061_), .Y(_12265_) );
	AOI21X1 AOI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_12021_), .B(_12066_), .C(_12265_), .Y(_12267_) );
	AOI21X1 AOI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_12261_), .B(_12262_), .C(_12260_), .Y(_12268_) );
	AOI21X1 AOI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_12258_), .B(_12253_), .C(_12218_), .Y(_12269_) );
	OAI21X1 OAI21X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_12268_), .B(_12269_), .C(_12267_), .Y(_12270_) );
	NAND3X1 NAND3X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_12270_), .B(_12264_), .C(_12191_), .Y(_12271_) );
	NAND3X1 NAND3X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_12186_), .B(_12180_), .C(_12184_), .Y(_12272_) );
	NAND3X1 NAND3X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_12147_), .B(_12188_), .C(_12187_), .Y(_12273_) );
	NAND2X1 NAND2X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_12272_), .B(_12273_), .Y(_12274_) );
	OAI21X1 OAI21X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_12268_), .B(_12269_), .C(_12193_), .Y(_12275_) );
	NAND3X1 NAND3X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_12259_), .B(_12263_), .C(_12267_), .Y(_12276_) );
	NAND3X1 NAND3X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_12275_), .B(_12276_), .C(_12274_), .Y(_12278_) );
	NAND3X1 NAND3X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_12271_), .B(_12278_), .C(_12145_), .Y(_12279_) );
	INVX1 INVX1_1775 ( .gnd(gnd), .vdd(vdd), .A(_12075_), .Y(_12280_) );
	AOI21X1 AOI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_12080_), .C(_12280_), .Y(_12281_) );
	AOI21X1 AOI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_12276_), .B(_12275_), .C(_12274_), .Y(_12282_) );
	AOI21X1 AOI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_12270_), .B(_12264_), .C(_12191_), .Y(_12283_) );
	OAI21X1 OAI21X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_12283_), .B(_12282_), .C(_12281_), .Y(_12284_) );
	NAND3X1 NAND3X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_12279_), .B(_12143_), .C(_12284_), .Y(_12285_) );
	NAND2X1 NAND2X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_12141_), .B(_12142_), .Y(_12286_) );
	OAI21X1 OAI21X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_12283_), .B(_12282_), .C(_12145_), .Y(_12287_) );
	NAND3X1 NAND3X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_12271_), .B(_12278_), .C(_12281_), .Y(_12289_) );
	NAND3X1 NAND3X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_12286_), .B(_12287_), .C(_12289_), .Y(_12290_) );
	NAND3X1 NAND3X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_12285_), .B(_12130_), .C(_12290_), .Y(_12291_) );
	AOI21X1 AOI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_11948_), .B(_12095_), .C(_12097_), .Y(_12292_) );
	AOI21X1 AOI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_12289_), .B(_12287_), .C(_12286_), .Y(_12293_) );
	AOI21X1 AOI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_12284_), .B(_12279_), .C(_12143_), .Y(_12294_) );
	OAI21X1 OAI21X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_12293_), .C(_12292_), .Y(_12295_) );
	NAND3X1 NAND3X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .B(_12291_), .C(_12295_), .Y(_12296_) );
	INVX1 INVX1_1776 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .Y(_12297_) );
	OAI21X1 OAI21X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_12293_), .C(_12130_), .Y(_12298_) );
	NAND3X1 NAND3X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_12285_), .B(_12290_), .C(_12292_), .Y(_12300_) );
	NAND3X1 NAND3X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .B(_12298_), .C(_12300_), .Y(_12301_) );
	AOI21X1 AOI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_12301_), .B(_12296_), .C(_12128_), .Y(_12302_) );
	NAND3X1 NAND3X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .B(_12291_), .C(_12295_), .Y(_12303_) );
	NAND3X1 NAND3X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .B(_12298_), .C(_12300_), .Y(_12304_) );
	AOI21X1 AOI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_12304_), .B(_12303_), .C(_12100_), .Y(_12305_) );
	AOI21X1 AOI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_11922_), .B(_11923_), .C(_17287_), .Y(_12306_) );
	AOI21X1 AOI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_12306_), .B(_12112_), .C(_12119_), .Y(_12307_) );
	OAI21X1 OAI21X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12305_), .C(_12307_), .Y(_12308_) );
	AOI21X1 AOI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_12301_), .B(_12296_), .C(_12100_), .Y(_12309_) );
	AOI21X1 AOI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_12304_), .B(_12303_), .C(_12128_), .Y(_12311_) );
	OAI21X1 OAI21X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_11928_), .B(_12121_), .C(_12109_), .Y(_12312_) );
	OAI21X1 OAI21X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .B(_12311_), .C(_12312_), .Y(_12313_) );
	NAND2X1 NAND2X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_12313_), .B(_12308_), .Y(_12314_) );
	XOR2X1 XOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_12127_), .B(_12314_), .Y(mulOut_15_) );
	AOI22X1 AOI22X1_281 ( .gnd(gnd), .vdd(vdd), .A(_12308_), .B(_12313_), .C(_12122_), .D(_12118_), .Y(_12315_) );
	INVX1 INVX1_1777 ( .gnd(gnd), .vdd(vdd), .A(_17303_), .Y(_12316_) );
	NAND2X1 NAND2X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_11933_), .B(_11927_), .Y(_12317_) );
	AOI22X1 AOI22X1_282 ( .gnd(gnd), .vdd(vdd), .A(_11935_), .B(_11925_), .C(_12317_), .D(_12316_), .Y(_12318_) );
	AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_12116_), .B(_12113_), .Y(_12319_) );
	NAND3X1 NAND3X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_12100_), .B(_12303_), .C(_12304_), .Y(_12321_) );
	NAND3X1 NAND3X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_12128_), .B(_12296_), .C(_12301_), .Y(_12322_) );
	AOI21X1 AOI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_12321_), .B(_12322_), .C(_12312_), .Y(_12323_) );
	NAND2X1 NAND2X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_12321_), .B(_12322_), .Y(_12324_) );
	NOR2X1 NOR2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_12307_), .B(_12324_), .Y(_12325_) );
	OAI22X1 OAI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(_12117_), .B(_12319_), .C(_12323_), .D(_12325_), .Y(_12326_) );
	NOR2X1 NOR2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_12125_), .B(_12113_), .Y(_12327_) );
	NOR2X1 NOR2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_11928_), .B(_12113_), .Y(_12328_) );
	AOI22X1 AOI22X1_283 ( .gnd(gnd), .vdd(vdd), .A(_12324_), .B(_12328_), .C(_12327_), .D(_12314_), .Y(_12329_) );
	OAI21X1 OAI21X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_12326_), .B(_12318_), .C(_12329_), .Y(_12330_) );
	AOI21X1 AOI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_11938_), .B(_12315_), .C(_12330_), .Y(_12331_) );
	OAI21X1 OAI21X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12305_), .C(_12119_), .Y(_12332_) );
	AOI21X1 AOI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_12290_), .B(_12285_), .C(_12130_), .Y(_12333_) );
	OAI21X1 OAI21X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_12129_), .B(_12333_), .C(_12291_), .Y(_12334_) );
	INVX1 INVX1_1778 ( .gnd(gnd), .vdd(vdd), .A(_12141_), .Y(_12335_) );
	AOI21X1 AOI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_12278_), .B(_12271_), .C(_12145_), .Y(_12336_) );
	OAI21X1 OAI21X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_12286_), .B(_12336_), .C(_12279_), .Y(_12337_) );
	NAND2X1 NAND2X1_2582 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf0), .B(adder_bOperand_16_bF_buf0), .Y(_12338_) );
	INVX1 INVX1_1779 ( .gnd(gnd), .vdd(vdd), .A(_12338_), .Y(_12339_) );
	NAND2X1 NAND2X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_12339_), .B(_12132_), .Y(_12340_) );
	INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_16_bF_buf3), .Y(_12342_) );
	NAND2X1 NAND2X1_2584 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf5), .B(adder_bOperand_15_bF_buf4), .Y(_12343_) );
	OAI21X1 OAI21X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf0), .B(_12342_), .C(_12343_), .Y(_12344_) );
	AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_12340_), .B(_12344_), .Y(_12345_) );
	OAI22X1 OAI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_11954_), .B(_12149_), .C(_12148_), .D(_12152_), .Y(_12346_) );
	NAND2X1 NAND2X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_12345_), .B(_12346_), .Y(_12347_) );
	INVX1 INVX1_1780 ( .gnd(gnd), .vdd(vdd), .A(_12347_), .Y(_12348_) );
	NOR2X1 NOR2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_12345_), .B(_12346_), .Y(_12349_) );
	NOR2X1 NOR2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_12349_), .B(_12348_), .Y(_12350_) );
	NOR2X1 NOR2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_12138_), .B(_12350_), .Y(_12351_) );
	NAND2X1 NAND2X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_12138_), .B(_12350_), .Y(_12354_) );
	INVX1 INVX1_1781 ( .gnd(gnd), .vdd(vdd), .A(_12354_), .Y(_12355_) );
	NOR2X1 NOR2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_12351_), .B(_12355_), .Y(_12356_) );
	NAND2X1 NAND2X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_12180_), .B(_12272_), .Y(_12357_) );
	NAND2X1 NAND2X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_12356_), .B(_12357_), .Y(_12358_) );
	OR2X2 OR2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_12357_), .B(_12356_), .Y(_12359_) );
	AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_12359_), .B(_12358_), .Y(_12360_) );
	AOI21X1 AOI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_12259_), .B(_12263_), .C(_12193_), .Y(_12361_) );
	OAI21X1 OAI21X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_12361_), .B(_12274_), .C(_12264_), .Y(_12362_) );
	NAND2X1 NAND2X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_12164_), .B(_12171_), .Y(_12363_) );
	INVX8 INVX8_71 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf1), .Y(_12365_) );
	NOR2X1 NOR2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf3), .B(_12365_), .Y(_12366_) );
	NAND2X1 NAND2X1_2590 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf1), .B(adder_bOperand_13_bF_buf1), .Y(_12367_) );
	OAI21X1 OAI21X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf2), .B(_17157_), .C(_12149_), .Y(_12368_) );
	OAI21X1 OAI21X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_12150_), .B(_12367_), .C(_12368_), .Y(_12369_) );
	XNOR2X1 XNOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_12369_), .B(_12366_), .Y(_12370_) );
	AOI22X1 AOI22X1_284 ( .gnd(gnd), .vdd(vdd), .A(_12166_), .B(_12167_), .C(_12156_), .D(_12160_), .Y(_12371_) );
	INVX1 INVX1_1782 ( .gnd(gnd), .vdd(vdd), .A(_12371_), .Y(_12372_) );
	NAND2X1 NAND2X1_2591 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf0), .B(adder_bOperand_11_bF_buf2), .Y(_12373_) );
	INVX1 INVX1_1783 ( .gnd(gnd), .vdd(vdd), .A(_12373_), .Y(_12374_) );
	NAND2X1 NAND2X1_2592 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf0), .B(adder_bOperand_9_bF_buf4), .Y(_12376_) );
	NOR2X1 NOR2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_12159_), .B(_12376_), .Y(_12377_) );
	INVX1 INVX1_1784 ( .gnd(gnd), .vdd(vdd), .A(_12377_), .Y(_12378_) );
	OAI21X1 OAI21X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_17025__bF_buf2), .C(_12159_), .Y(_12379_) );
	NAND3X1 NAND3X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_12374_), .B(_12379_), .C(_12378_), .Y(_12380_) );
	AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_12159_), .B(_12376_), .Y(_12381_) );
	OAI21X1 OAI21X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_12377_), .B(_12381_), .C(_12373_), .Y(_12382_) );
	NAND3X1 NAND3X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_12382_), .B(_12380_), .C(_12372_), .Y(_12383_) );
	NOR3X1 NOR3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_12373_), .B(_12377_), .C(_12381_), .Y(_12384_) );
	AOI22X1 AOI22X1_285 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf4), .B(adder_bOperand_11_bF_buf1), .C(_12379_), .D(_12378_), .Y(_12385_) );
	OAI21X1 OAI21X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_12384_), .B(_12385_), .C(_12371_), .Y(_12387_) );
	NAND3X1 NAND3X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_12383_), .C(_12387_), .Y(_12388_) );
	INVX1 INVX1_1785 ( .gnd(gnd), .vdd(vdd), .A(_12366_), .Y(_12389_) );
	OR2X2 OR2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_12369_), .B(_12389_), .Y(_12390_) );
	OAI21X1 OAI21X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf2), .B(_12365_), .C(_12369_), .Y(_12391_) );
	NAND2X1 NAND2X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_12391_), .B(_12390_), .Y(_12392_) );
	OAI21X1 OAI21X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_12384_), .B(_12385_), .C(_12372_), .Y(_12393_) );
	NAND3X1 NAND3X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_12371_), .B(_12382_), .C(_12380_), .Y(_12394_) );
	NAND3X1 NAND3X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_12394_), .B(_12392_), .C(_12393_), .Y(_12395_) );
	AOI21X1 AOI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_12199_), .B(_12200_), .C(_12205_), .Y(_12396_) );
	OAI21X1 OAI21X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_12214_), .B(_12396_), .C(_12206_), .Y(_12398_) );
	AOI21X1 AOI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_12388_), .B(_12395_), .C(_12398_), .Y(_12399_) );
	AOI21X1 AOI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_12393_), .B(_12394_), .C(_12392_), .Y(_12400_) );
	AOI22X1 AOI22X1_286 ( .gnd(gnd), .vdd(vdd), .A(_12390_), .B(_12391_), .C(_12383_), .D(_12387_), .Y(_12401_) );
	NOR3X1 NOR3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_12204_), .B(_12210_), .C(_12207_), .Y(_12402_) );
	AOI21X1 AOI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_12211_), .B(_12194_), .C(_12402_), .Y(_12403_) );
	NOR3X1 NOR3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_12401_), .B(_12400_), .C(_12403_), .Y(_12404_) );
	OAI21X1 OAI21X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_12399_), .B(_12404_), .C(_12363_), .Y(_12405_) );
	AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_12171_), .B(_12164_), .Y(_12406_) );
	OAI21X1 OAI21X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_12401_), .B(_12400_), .C(_12403_), .Y(_12407_) );
	NAND3X1 NAND3X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_12388_), .B(_12395_), .C(_12398_), .Y(_12409_) );
	NAND3X1 NAND3X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_12406_), .B(_12407_), .C(_12409_), .Y(_12410_) );
	NAND2X1 NAND2X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_12410_), .B(_12405_), .Y(_12411_) );
	AOI21X1 AOI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_12248_), .B(_12252_), .C(_12219_), .Y(_12412_) );
	OAI21X1 OAI21X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_12412_), .B(_12260_), .C(_12253_), .Y(_12413_) );
	OAI21X1 OAI21X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_12195_), .B(_12198_), .C(_12209_), .Y(_12414_) );
	NOR2X1 NOR2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_14728__bF_buf2), .Y(_12415_) );
	NAND2X1 NAND2X1_2595 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf3), .B(aOperand_frameOut_10_bF_buf3), .Y(_12416_) );
	INVX1 INVX1_1786 ( .gnd(gnd), .vdd(vdd), .A(_12416_), .Y(_12417_) );
	NAND2X1 NAND2X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_12208_), .B(_12417_), .Y(_12418_) );
	OAI21X1 OAI21X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf0), .B(_16940_), .C(_12196_), .Y(_12420_) );
	NAND3X1 NAND3X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_12415_), .B(_12420_), .C(_12418_), .Y(_12421_) );
	INVX1 INVX1_1787 ( .gnd(gnd), .vdd(vdd), .A(_12415_), .Y(_12422_) );
	OAI21X1 OAI21X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_13830_), .B(_15812__bF_buf0), .C(_12417_), .Y(_12423_) );
	OAI21X1 OAI21X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf3), .B(_16940_), .C(_12208_), .Y(_12424_) );
	NAND3X1 NAND3X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_12423_), .B(_12422_), .C(_12424_), .Y(_12425_) );
	NOR2X1 NOR2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_12202_), .B(_12222_), .Y(_12426_) );
	AOI21X1 AOI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_12224_), .B(_12221_), .C(_12426_), .Y(_12427_) );
	INVX1 INVX1_1788 ( .gnd(gnd), .vdd(vdd), .A(_12427_), .Y(_12428_) );
	NAND3X1 NAND3X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_12421_), .B(_12425_), .C(_12428_), .Y(_12429_) );
	AOI21X1 AOI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_12423_), .B(_12424_), .C(_12422_), .Y(_12431_) );
	AOI21X1 AOI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_12418_), .B(_12420_), .C(_12415_), .Y(_12432_) );
	OAI21X1 OAI21X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_12432_), .B(_12431_), .C(_12427_), .Y(_12433_) );
	NAND3X1 NAND3X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_12414_), .B(_12429_), .C(_12433_), .Y(_12434_) );
	INVX1 INVX1_1789 ( .gnd(gnd), .vdd(vdd), .A(_12414_), .Y(_12435_) );
	NAND3X1 NAND3X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_12421_), .B(_12427_), .C(_12425_), .Y(_12436_) );
	OAI21X1 OAI21X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_12432_), .B(_12431_), .C(_12428_), .Y(_12437_) );
	NAND3X1 NAND3X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_12436_), .B(_12435_), .C(_12437_), .Y(_12438_) );
	AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_12434_), .B(_12438_), .Y(_12439_) );
	AOI21X1 AOI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_12235_), .B(_12239_), .C(_12227_), .Y(_12440_) );
	OAI21X1 OAI21X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_12440_), .B(_12249_), .C(_12240_), .Y(_12442_) );
	NAND2X1 NAND2X1_2597 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf4), .B(aOperand_frameOut_11_bF_buf2), .Y(_12443_) );
	INVX1 INVX1_1790 ( .gnd(gnd), .vdd(vdd), .A(_12443_), .Y(_12444_) );
	AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf3), .B(aOperand_frameOut_12_bF_buf0), .Y(_12445_) );
	AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf3), .B(aOperand_frameOut_13_bF_buf0), .Y(_12446_) );
	NAND2X1 NAND2X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_12445_), .B(_12446_), .Y(_12447_) );
	OAI21X1 OAI21X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf0), .B(_11858_), .C(_12222_), .Y(_12448_) );
	NAND3X1 NAND3X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_12444_), .B(_12448_), .C(_12447_), .Y(_12449_) );
	OAI21X1 OAI21X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_17236__bF_buf3), .C(_12446_), .Y(_12450_) );
	OAI21X1 OAI21X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf3), .B(_11858_), .C(_12445_), .Y(_12451_) );
	NAND3X1 NAND3X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_12443_), .B(_12450_), .C(_12451_), .Y(_12453_) );
	AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_12453_), .B(_12449_), .Y(_12454_) );
	OAI21X1 OAI21X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_12228_), .B(_12238_), .C(_12232_), .Y(_12455_) );
	NAND2X1 NAND2X1_2599 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf2), .B(aOperand_frameOut_14_bF_buf2), .Y(_12456_) );
	INVX1 INVX1_1791 ( .gnd(gnd), .vdd(vdd), .A(_12456_), .Y(_12457_) );
	AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf3), .B(aOperand_frameOut_15_bF_buf3), .Y(_12458_) );
	AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(aOperand_frameOut_16_bF_buf0), .Y(_12459_) );
	NAND2X1 NAND2X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_12458_), .B(_12459_), .Y(_12460_) );
	INVX4 INVX4_17 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_16_bF_buf4), .Y(_12461_) );
	OAI22X1 OAI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf1), .B(_12461_), .C(_11776__bF_buf0), .D(_12233_), .Y(_12462_) );
	NAND3X1 NAND3X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_12457_), .B(_12462_), .C(_12460_), .Y(_12464_) );
	NAND2X1 NAND2X1_2601 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .B(aOperand_frameOut_16_bF_buf3), .Y(_12465_) );
	NOR2X1 NOR2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_12236_), .B(_12465_), .Y(_12466_) );
	AOI21X1 AOI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .B(aOperand_frameOut_16_bF_buf2), .C(_12458_), .Y(_12467_) );
	OAI21X1 OAI21X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_12466_), .B(_12467_), .C(_12456_), .Y(_12468_) );
	NAND3X1 NAND3X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_12464_), .B(_12455_), .C(_12468_), .Y(_12469_) );
	AOI21X1 AOI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_12234_), .B(_12229_), .C(_12237_), .Y(_12470_) );
	OAI21X1 OAI21X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf3), .B(_12233_), .C(_12459_), .Y(_12471_) );
	OAI21X1 OAI21X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf0), .B(_12461_), .C(_12458_), .Y(_12472_) );
	AOI21X1 AOI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_12471_), .B(_12472_), .C(_12456_), .Y(_12473_) );
	AOI21X1 AOI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_12460_), .B(_12462_), .C(_12457_), .Y(_12475_) );
	OAI21X1 OAI21X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_12475_), .B(_12473_), .C(_12470_), .Y(_12476_) );
	NAND3X1 NAND3X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_12454_), .B(_12469_), .C(_12476_), .Y(_12477_) );
	NAND2X1 NAND2X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_12449_), .B(_12453_), .Y(_12478_) );
	OAI21X1 OAI21X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_12475_), .B(_12473_), .C(_12455_), .Y(_12479_) );
	NAND3X1 NAND3X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_12464_), .B(_12470_), .C(_12468_), .Y(_12480_) );
	NAND3X1 NAND3X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_12478_), .B(_12480_), .C(_12479_), .Y(_12481_) );
	NAND3X1 NAND3X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_12477_), .B(_12481_), .C(_12442_), .Y(_12482_) );
	INVX1 INVX1_1792 ( .gnd(gnd), .vdd(vdd), .A(_12240_), .Y(_12483_) );
	AOI21X1 AOI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_12226_), .B(_12247_), .C(_12483_), .Y(_12484_) );
	AOI21X1 AOI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_12479_), .B(_12480_), .C(_12478_), .Y(_12486_) );
	AOI21X1 AOI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_12476_), .B(_12469_), .C(_12454_), .Y(_12487_) );
	OAI21X1 OAI21X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_12486_), .B(_12487_), .C(_12484_), .Y(_12488_) );
	NAND3X1 NAND3X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_12482_), .B(_12439_), .C(_12488_), .Y(_12489_) );
	NAND2X1 NAND2X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_12438_), .B(_12434_), .Y(_12490_) );
	NAND2X1 NAND2X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_12477_), .B(_12481_), .Y(_12491_) );
	NOR2X1 NOR2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_12484_), .B(_12491_), .Y(_12492_) );
	AOI21X1 AOI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_12477_), .B(_12481_), .C(_12442_), .Y(_12493_) );
	OAI21X1 OAI21X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_12493_), .B(_12492_), .C(_12490_), .Y(_12494_) );
	NAND3X1 NAND3X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_12413_), .B(_12489_), .C(_12494_), .Y(_12495_) );
	NAND2X1 NAND2X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_12248_), .B(_12252_), .Y(_12497_) );
	NOR2X1 NOR2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_12254_), .B(_12497_), .Y(_12498_) );
	AOI21X1 AOI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_12218_), .B(_12258_), .C(_12498_), .Y(_12499_) );
	OAI21X1 OAI21X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_12486_), .B(_12487_), .C(_12442_), .Y(_12500_) );
	NAND3X1 NAND3X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_12477_), .B(_12481_), .C(_12484_), .Y(_12501_) );
	AOI21X1 AOI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_12501_), .B(_12500_), .C(_12490_), .Y(_12502_) );
	AOI21X1 AOI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_12488_), .B(_12482_), .C(_12439_), .Y(_12503_) );
	OAI21X1 OAI21X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_12503_), .B(_12502_), .C(_12499_), .Y(_12504_) );
	NAND3X1 NAND3X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_12495_), .B(_12504_), .C(_12411_), .Y(_12505_) );
	NAND3X1 NAND3X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .B(_12407_), .C(_12409_), .Y(_12506_) );
	OAI21X1 OAI21X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_12399_), .B(_12404_), .C(_12406_), .Y(_12508_) );
	NAND2X1 NAND2X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_12506_), .B(_12508_), .Y(_12509_) );
	OAI21X1 OAI21X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_12503_), .B(_12502_), .C(_12413_), .Y(_12510_) );
	NAND3X1 NAND3X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_12489_), .B(_12494_), .C(_12499_), .Y(_12511_) );
	NAND3X1 NAND3X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_12510_), .B(_12511_), .C(_12509_), .Y(_12512_) );
	NAND3X1 NAND3X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_12505_), .B(_12512_), .C(_12362_), .Y(_12513_) );
	INVX1 INVX1_1793 ( .gnd(gnd), .vdd(vdd), .A(_12264_), .Y(_12514_) );
	AOI21X1 AOI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_12191_), .B(_12270_), .C(_12514_), .Y(_12515_) );
	AOI21X1 AOI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_12511_), .B(_12510_), .C(_12509_), .Y(_12516_) );
	AOI21X1 AOI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_12495_), .B(_12504_), .C(_12411_), .Y(_12517_) );
	OAI21X1 OAI21X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_12517_), .B(_12516_), .C(_12515_), .Y(_12519_) );
	NAND3X1 NAND3X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_12513_), .B(_12519_), .C(_12360_), .Y(_12520_) );
	NAND2X1 NAND2X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12359_), .Y(_12521_) );
	OAI21X1 OAI21X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_12517_), .B(_12516_), .C(_12362_), .Y(_12522_) );
	NAND3X1 NAND3X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_12505_), .B(_12512_), .C(_12515_), .Y(_12523_) );
	NAND3X1 NAND3X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_12521_), .B(_12522_), .C(_12523_), .Y(_12524_) );
	NAND3X1 NAND3X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_12337_), .B(_12520_), .C(_12524_), .Y(_12525_) );
	INVX1 INVX1_1794 ( .gnd(gnd), .vdd(vdd), .A(_12279_), .Y(_12526_) );
	AOI21X1 AOI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_12143_), .B(_12284_), .C(_12526_), .Y(_12527_) );
	AOI21X1 AOI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_12523_), .B(_12522_), .C(_12521_), .Y(_12528_) );
	AOI21X1 AOI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_12519_), .B(_12513_), .C(_12360_), .Y(_12530_) );
	OAI21X1 OAI21X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_12530_), .B(_12528_), .C(_12527_), .Y(_12531_) );
	NAND3X1 NAND3X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_12335_), .B(_12525_), .C(_12531_), .Y(_12532_) );
	OAI21X1 OAI21X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_12530_), .B(_12528_), .C(_12337_), .Y(_12533_) );
	NAND3X1 NAND3X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_12520_), .B(_12524_), .C(_12527_), .Y(_12534_) );
	NAND3X1 NAND3X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_12141_), .B(_12533_), .C(_12534_), .Y(_12535_) );
	NAND3X1 NAND3X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_12532_), .B(_12535_), .C(_12334_), .Y(_12536_) );
	INVX1 INVX1_1795 ( .gnd(gnd), .vdd(vdd), .A(_12291_), .Y(_12537_) );
	AOI21X1 AOI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .B(_12295_), .C(_12537_), .Y(_12538_) );
	AOI21X1 AOI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_12534_), .B(_12533_), .C(_12141_), .Y(_12539_) );
	AOI21X1 AOI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_12531_), .B(_12525_), .C(_12335_), .Y(_12541_) );
	OAI21X1 OAI21X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_12541_), .B(_12539_), .C(_12538_), .Y(_12542_) );
	NAND3X1 NAND3X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_12536_), .B(_12309_), .C(_12542_), .Y(_12543_) );
	NAND3X1 NAND3X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_12128_), .B(_12303_), .C(_12304_), .Y(_12544_) );
	OAI21X1 OAI21X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_12541_), .B(_12539_), .C(_12334_), .Y(_12545_) );
	NAND3X1 NAND3X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_12532_), .B(_12535_), .C(_12538_), .Y(_12546_) );
	NAND3X1 NAND3X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_12544_), .B(_12545_), .C(_12546_), .Y(_12547_) );
	NAND3X1 NAND3X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_12543_), .B(_12547_), .C(_12332_), .Y(_12548_) );
	AOI21X1 AOI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_12322_), .B(_12321_), .C(_12109_), .Y(_12549_) );
	NAND3X1 NAND3X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_12544_), .B(_12536_), .C(_12542_), .Y(_12550_) );
	NAND3X1 NAND3X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .B(_12545_), .C(_12546_), .Y(_12552_) );
	NAND3X1 NAND3X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_12549_), .B(_12550_), .C(_12552_), .Y(_12553_) );
	NAND2X1 NAND2X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_12553_), .B(_12548_), .Y(_12554_) );
	XNOR2X1 XNOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_12331_), .B(_12554_), .Y(mulOut_16_) );
	INVX1 INVX1_1796 ( .gnd(gnd), .vdd(vdd), .A(_12331_), .Y(_12555_) );
	AOI21X1 AOI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_12552_), .B(_12550_), .C(_12332_), .Y(_12556_) );
	AOI21X1 AOI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_12555_), .B(_12554_), .C(_12556_), .Y(_12557_) );
	INVX1 INVX1_1797 ( .gnd(gnd), .vdd(vdd), .A(_12536_), .Y(_12558_) );
	AOI21X1 AOI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_12524_), .B(_12520_), .C(_12337_), .Y(_12559_) );
	OAI21X1 OAI21X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_12141_), .B(_12559_), .C(_12525_), .Y(_12560_) );
	INVX1 INVX1_1798 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .Y(_12562_) );
	AOI21X1 AOI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_12505_), .B(_12512_), .C(_12362_), .Y(_12563_) );
	OAI21X1 OAI21X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_12521_), .B(_12563_), .C(_12513_), .Y(_12564_) );
	OAI21X1 OAI21X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_12406_), .B(_12399_), .C(_12409_), .Y(_12565_) );
	INVX4 INVX4_18 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_17_bF_buf0), .Y(_12566_) );
	NOR2X1 NOR2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf3), .B(_12566_), .Y(_12567_) );
	NAND2X1 NAND2X1_2609 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf4), .B(adder_bOperand_15_bF_buf3), .Y(_12568_) );
	INVX1 INVX1_1799 ( .gnd(gnd), .vdd(vdd), .A(_12568_), .Y(_12569_) );
	NAND2X1 NAND2X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_12339_), .B(_12569_), .Y(_12570_) );
	OAI21X1 OAI21X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf1), .B(_12131_), .C(_12338_), .Y(_12571_) );
	NAND3X1 NAND3X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_12567_), .B(_12571_), .C(_12570_), .Y(_12573_) );
	NAND2X1 NAND2X1_2611 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf3), .B(adder_bOperand_16_bF_buf2), .Y(_12574_) );
	OAI21X1 OAI21X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_12343_), .B(_12574_), .C(_12571_), .Y(_12575_) );
	OAI21X1 OAI21X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf2), .B(_12566_), .C(_12575_), .Y(_12576_) );
	NAND2X1 NAND2X1_2612 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf0), .B(adder_bOperand_12_bF_buf3), .Y(_12577_) );
	NOR2X1 NOR2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_12149_), .B(_12577_), .Y(_12578_) );
	AOI21X1 AOI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_12368_), .B(_12366_), .C(_12578_), .Y(_12579_) );
	INVX1 INVX1_1800 ( .gnd(gnd), .vdd(vdd), .A(_12579_), .Y(_12580_) );
	NAND3X1 NAND3X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_12573_), .B(_12576_), .C(_12580_), .Y(_12581_) );
	AOI21X1 AOI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_12576_), .B(_12573_), .C(_12580_), .Y(_12582_) );
	INVX1 INVX1_1801 ( .gnd(gnd), .vdd(vdd), .A(_12582_), .Y(_12583_) );
	NAND2X1 NAND2X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_12583_), .Y(_12584_) );
	NAND2X1 NAND2X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_12340_), .B(_12347_), .Y(_12585_) );
	XNOR2X1 XNOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_12584_), .B(_12585_), .Y(_12586_) );
	NAND2X1 NAND2X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_12586_), .B(_12565_), .Y(_12587_) );
	AOI21X1 AOI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_12363_), .B(_12407_), .C(_12404_), .Y(_12588_) );
	XOR2X1 XOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_12584_), .B(_12585_), .Y(_12589_) );
	NAND2X1 NAND2X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_12589_), .B(_12588_), .Y(_12590_) );
	NAND3X1 NAND3X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_12354_), .B(_12587_), .C(_12590_), .Y(_12591_) );
	NAND2X1 NAND2X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_12586_), .B(_12588_), .Y(_12592_) );
	NAND2X1 NAND2X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_12589_), .B(_12565_), .Y(_12594_) );
	NAND3X1 NAND3X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_12355_), .B(_12594_), .C(_12592_), .Y(_12595_) );
	NAND2X1 NAND2X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_12591_), .B(_12595_), .Y(_12596_) );
	AOI21X1 AOI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_12494_), .B(_12489_), .C(_12413_), .Y(_12597_) );
	OAI21X1 OAI21X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_12509_), .B(_12597_), .C(_12495_), .Y(_12598_) );
	NAND2X1 NAND2X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_12383_), .B(_12388_), .Y(_12599_) );
	NAND2X1 NAND2X1_2621 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf3), .B(adder_bOperand_14_bF_buf0), .Y(_12600_) );
	INVX1 INVX1_1802 ( .gnd(gnd), .vdd(vdd), .A(_12600_), .Y(_12601_) );
	NAND2X1 NAND2X1_2622 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf3), .B(adder_bOperand_13_bF_buf0), .Y(_12602_) );
	OAI21X1 OAI21X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_17157_), .C(_12367_), .Y(_12603_) );
	OAI21X1 OAI21X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_12577_), .B(_12602_), .C(_12603_), .Y(_12604_) );
	XNOR2X1 XNOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_12604_), .B(_12601_), .Y(_12605_) );
	OAI21X1 OAI21X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_12373_), .B(_12381_), .C(_12378_), .Y(_12606_) );
	NAND2X1 NAND2X1_2623 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf0), .B(adder_bOperand_11_bF_buf0), .Y(_12607_) );
	INVX1 INVX1_1803 ( .gnd(gnd), .vdd(vdd), .A(_12607_), .Y(_12608_) );
	AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf4), .B(adder_bOperand_10_bF_buf2), .Y(_12609_) );
	AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf2), .B(adder_bOperand_9_bF_buf3), .Y(_12610_) );
	NAND2X1 NAND2X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_12609_), .B(_12610_), .Y(_12611_) );
	OAI22X1 OAI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_16887_), .C(_15035_), .D(_17025__bF_buf1), .Y(_12612_) );
	NAND3X1 NAND3X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_12608_), .B(_12612_), .C(_12611_), .Y(_12613_) );
	OAI21X1 OAI21X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_16887_), .C(_12610_), .Y(_12616_) );
	OAI21X1 OAI21X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_17025__bF_buf0), .C(_12609_), .Y(_12617_) );
	NAND3X1 NAND3X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_12607_), .B(_12616_), .C(_12617_), .Y(_12618_) );
	NAND3X1 NAND3X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_12613_), .B(_12618_), .C(_12606_), .Y(_12619_) );
	AOI21X1 AOI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_12379_), .B(_12374_), .C(_12377_), .Y(_12620_) );
	AOI21X1 AOI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_12616_), .B(_12617_), .C(_12607_), .Y(_12621_) );
	AOI21X1 AOI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_12611_), .B(_12612_), .C(_12608_), .Y(_12622_) );
	OAI21X1 OAI21X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_12622_), .B(_12621_), .C(_12620_), .Y(_12623_) );
	NAND3X1 NAND3X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_12623_), .B(_12619_), .C(_12605_), .Y(_12624_) );
	XNOR2X1 XNOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_12604_), .B(_12600_), .Y(_12625_) );
	OAI21X1 OAI21X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_12622_), .B(_12621_), .C(_12606_), .Y(_12627_) );
	NAND3X1 NAND3X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_12613_), .B(_12620_), .C(_12618_), .Y(_12628_) );
	NAND3X1 NAND3X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_12627_), .B(_12628_), .C(_12625_), .Y(_12629_) );
	AOI21X1 AOI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_12421_), .B(_12425_), .C(_12428_), .Y(_12630_) );
	OAI21X1 OAI21X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_12435_), .B(_12630_), .C(_12429_), .Y(_12631_) );
	AOI21X1 AOI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_12624_), .B(_12629_), .C(_12631_), .Y(_12632_) );
	NAND2X1 NAND2X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_12624_), .B(_12629_), .Y(_12633_) );
	NAND2X1 NAND2X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_12421_), .B(_12425_), .Y(_12634_) );
	NOR2X1 NOR2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_12427_), .B(_12634_), .Y(_12635_) );
	AOI21X1 AOI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_12433_), .B(_12414_), .C(_12635_), .Y(_12636_) );
	NOR2X1 NOR2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_12636_), .B(_12633_), .Y(_12638_) );
	OAI21X1 OAI21X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_12632_), .B(_12638_), .C(_12599_), .Y(_12639_) );
	INVX1 INVX1_1804 ( .gnd(gnd), .vdd(vdd), .A(_12599_), .Y(_12640_) );
	NAND2X1 NAND2X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_12636_), .B(_12633_), .Y(_12641_) );
	NAND3X1 NAND3X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_12624_), .B(_12629_), .C(_12631_), .Y(_12642_) );
	NAND3X1 NAND3X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_12642_), .B(_12641_), .C(_12640_), .Y(_12643_) );
	NAND2X1 NAND2X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_12643_), .B(_12639_), .Y(_12644_) );
	OAI21X1 OAI21X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_12490_), .B(_12493_), .C(_12482_), .Y(_12645_) );
	AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_12421_), .B(_12418_), .Y(_12646_) );
	NOR2X1 NOR2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf1), .B(_15812__bF_buf3), .Y(_12647_) );
	AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf3), .B(aOperand_frameOut_11_bF_buf1), .Y(_12649_) );
	NAND2X1 NAND2X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_12649_), .B(_12417_), .Y(_12650_) );
	NAND2X1 NAND2X1_2630 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf2), .B(aOperand_frameOut_10_bF_buf2), .Y(_12651_) );
	OAI21X1 OAI21X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf2), .B(_17077_), .C(_12651_), .Y(_12652_) );
	NAND3X1 NAND3X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_12647_), .B(_12652_), .C(_12650_), .Y(_12653_) );
	INVX1 INVX1_1805 ( .gnd(gnd), .vdd(vdd), .A(_12647_), .Y(_12654_) );
	NAND3X1 NAND3X1_2690 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf2), .B(aOperand_frameOut_11_bF_buf0), .C(_12651_), .Y(_12655_) );
	NAND2X1 NAND2X1_2631 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf1), .B(aOperand_frameOut_11_bF_buf4), .Y(_12656_) );
	NAND3X1 NAND3X1_2691 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf1), .B(aOperand_frameOut_10_bF_buf1), .C(_12656_), .Y(_12657_) );
	NAND3X1 NAND3X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_12655_), .B(_12657_), .C(_12654_), .Y(_12658_) );
	NAND2X1 NAND2X1_2632 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf2), .B(aOperand_frameOut_13_bF_buf4), .Y(_12660_) );
	NOR2X1 NOR2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_12222_), .B(_12660_), .Y(_12661_) );
	AOI21X1 AOI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_12448_), .B(_12444_), .C(_12661_), .Y(_12662_) );
	INVX1 INVX1_1806 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .Y(_12663_) );
	NAND3X1 NAND3X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_12653_), .B(_12658_), .C(_12663_), .Y(_12664_) );
	AOI21X1 AOI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_12655_), .B(_12657_), .C(_12654_), .Y(_12665_) );
	AOI21X1 AOI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_12650_), .B(_12652_), .C(_12647_), .Y(_12666_) );
	OAI21X1 OAI21X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_12665_), .B(_12666_), .C(_12662_), .Y(_12667_) );
	NAND3X1 NAND3X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_12646_), .B(_12667_), .C(_12664_), .Y(_12668_) );
	OAI21X1 OAI21X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_12196_), .B(_12416_), .C(_12421_), .Y(_12669_) );
	NAND3X1 NAND3X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .B(_12653_), .C(_12658_), .Y(_12671_) );
	OAI21X1 OAI21X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_12665_), .B(_12666_), .C(_12663_), .Y(_12672_) );
	NAND3X1 NAND3X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_12669_), .B(_12671_), .C(_12672_), .Y(_12673_) );
	NAND2X1 NAND2X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_12673_), .B(_12668_), .Y(_12674_) );
	AOI21X1 AOI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_12468_), .B(_12464_), .C(_12455_), .Y(_12675_) );
	OAI21X1 OAI21X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_12478_), .B(_12675_), .C(_12469_), .Y(_12676_) );
	NAND2X1 NAND2X1_2634 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf3), .B(aOperand_frameOut_12_bF_buf4), .Y(_12677_) );
	AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf2), .B(aOperand_frameOut_13_bF_buf3), .Y(_12678_) );
	AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf1), .B(aOperand_frameOut_14_bF_buf1), .Y(_12679_) );
	NAND2X1 NAND2X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_12678_), .B(_12679_), .Y(_12680_) );
	NAND2X1 NAND2X1_2636 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf1), .B(aOperand_frameOut_13_bF_buf2), .Y(_12682_) );
	OAI21X1 OAI21X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf2), .B(_12039_), .C(_12682_), .Y(_12683_) );
	NAND3X1 NAND3X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_12677_), .B(_12683_), .C(_12680_), .Y(_12684_) );
	INVX1 INVX1_1807 ( .gnd(gnd), .vdd(vdd), .A(_12677_), .Y(_12685_) );
	NAND2X1 NAND2X1_2637 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf0), .B(aOperand_frameOut_14_bF_buf0), .Y(_12686_) );
	NOR2X1 NOR2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_12660_), .B(_12686_), .Y(_12687_) );
	NOR2X1 NOR2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_12678_), .B(_12679_), .Y(_12688_) );
	OAI21X1 OAI21X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_12687_), .B(_12688_), .C(_12685_), .Y(_12689_) );
	NAND2X1 NAND2X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_12684_), .B(_12689_), .Y(_12690_) );
	OAI21X1 OAI21X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_12456_), .B(_12467_), .C(_12460_), .Y(_12691_) );
	NAND2X1 NAND2X1_2639 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf1), .B(aOperand_frameOut_15_bF_buf2), .Y(_12693_) );
	INVX1 INVX1_1808 ( .gnd(gnd), .vdd(vdd), .A(_12693_), .Y(_12694_) );
	AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf1), .B(aOperand_frameOut_16_bF_buf1), .Y(_12695_) );
	AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(aOperand_frameOut_17_bF_buf1), .Y(_12696_) );
	NAND2X1 NAND2X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_12695_), .B(_12696_), .Y(_12697_) );
	NAND2X1 NAND2X1_2641 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .B(aOperand_frameOut_17_bF_buf0), .Y(_12698_) );
	NAND2X1 NAND2X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12698_), .Y(_12699_) );
	NAND3X1 NAND3X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_12694_), .B(_12699_), .C(_12697_), .Y(_12700_) );
	NOR2X1 NOR2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12698_), .Y(_12701_) );
	AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_12465_), .B(_12698_), .Y(_12702_) );
	OAI21X1 OAI21X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_12701_), .B(_12702_), .C(_12693_), .Y(_12704_) );
	NAND3X1 NAND3X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_12700_), .B(_12704_), .C(_12691_), .Y(_12705_) );
	AOI21X1 AOI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_12462_), .B(_12457_), .C(_12466_), .Y(_12706_) );
	OAI21X1 OAI21X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf2), .B(_12461_), .C(_12696_), .Y(_12707_) );
	INVX4 INVX4_19 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_17_bF_buf4), .Y(_12708_) );
	OAI21X1 OAI21X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf4), .B(_12708_), .C(_12695_), .Y(_12709_) );
	AOI21X1 AOI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_12707_), .B(_12709_), .C(_12693_), .Y(_12710_) );
	AOI21X1 AOI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_12697_), .B(_12699_), .C(_12694_), .Y(_12711_) );
	OAI21X1 OAI21X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_12711_), .B(_12710_), .C(_12706_), .Y(_12712_) );
	NAND3X1 NAND3X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_12690_), .B(_12705_), .C(_12712_), .Y(_12713_) );
	NAND3X1 NAND3X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_12685_), .B(_12683_), .C(_12680_), .Y(_12715_) );
	OAI21X1 OAI21X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_12687_), .B(_12688_), .C(_12677_), .Y(_12716_) );
	NAND2X1 NAND2X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_12715_), .B(_12716_), .Y(_12717_) );
	OAI21X1 OAI21X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_12711_), .B(_12710_), .C(_12691_), .Y(_12718_) );
	NAND3X1 NAND3X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_12700_), .B(_12706_), .C(_12704_), .Y(_12719_) );
	NAND3X1 NAND3X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_12717_), .B(_12719_), .C(_12718_), .Y(_12720_) );
	NAND3X1 NAND3X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_12720_), .B(_12713_), .C(_12676_), .Y(_12721_) );
	NOR3X1 NOR3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_12470_), .B(_12475_), .C(_12473_), .Y(_12722_) );
	AOI21X1 AOI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_12454_), .B(_12476_), .C(_12722_), .Y(_12723_) );
	AOI21X1 AOI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_12718_), .B(_12719_), .C(_12717_), .Y(_12724_) );
	AOI21X1 AOI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_12712_), .B(_12705_), .C(_12690_), .Y(_12726_) );
	OAI21X1 OAI21X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_12724_), .B(_12726_), .C(_12723_), .Y(_12727_) );
	NAND3X1 NAND3X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_12721_), .B(_12674_), .C(_12727_), .Y(_12728_) );
	NAND3X1 NAND3X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_12669_), .B(_12667_), .C(_12664_), .Y(_12729_) );
	NAND3X1 NAND3X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_12646_), .B(_12671_), .C(_12672_), .Y(_12730_) );
	NAND2X1 NAND2X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_12730_), .B(_12729_), .Y(_12731_) );
	OAI21X1 OAI21X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_12724_), .B(_12726_), .C(_12676_), .Y(_12732_) );
	NAND3X1 NAND3X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_12713_), .B(_12720_), .C(_12723_), .Y(_12733_) );
	NAND3X1 NAND3X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_12731_), .B(_12733_), .C(_12732_), .Y(_12734_) );
	NAND3X1 NAND3X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_12728_), .B(_12734_), .C(_12645_), .Y(_12735_) );
	AOI21X1 AOI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_12439_), .B(_12488_), .C(_12492_), .Y(_12737_) );
	AOI21X1 AOI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_12732_), .B(_12733_), .C(_12731_), .Y(_12738_) );
	AOI21X1 AOI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_12727_), .B(_12721_), .C(_12674_), .Y(_12739_) );
	OAI21X1 OAI21X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_12738_), .B(_12739_), .C(_12737_), .Y(_12740_) );
	NAND3X1 NAND3X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_12735_), .B(_12740_), .C(_12644_), .Y(_12741_) );
	NAND3X1 NAND3X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_12599_), .B(_12642_), .C(_12641_), .Y(_12742_) );
	OAI21X1 OAI21X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_12632_), .B(_12638_), .C(_12640_), .Y(_12743_) );
	NAND2X1 NAND2X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_12742_), .B(_12743_), .Y(_12744_) );
	OAI21X1 OAI21X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_12738_), .B(_12739_), .C(_12645_), .Y(_12745_) );
	NAND3X1 NAND3X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_12728_), .B(_12734_), .C(_12737_), .Y(_12746_) );
	NAND3X1 NAND3X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_12745_), .B(_12746_), .C(_12744_), .Y(_12748_) );
	NAND3X1 NAND3X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_12741_), .B(_12748_), .C(_12598_), .Y(_12749_) );
	NOR3X1 NOR3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_12503_), .B(_12502_), .C(_12499_), .Y(_12750_) );
	AOI21X1 AOI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_12411_), .B(_12504_), .C(_12750_), .Y(_12751_) );
	AOI21X1 AOI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_12746_), .B(_12745_), .C(_12744_), .Y(_12752_) );
	AOI21X1 AOI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_12740_), .B(_12735_), .C(_12644_), .Y(_12753_) );
	OAI21X1 OAI21X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_12752_), .B(_12753_), .C(_12751_), .Y(_12754_) );
	NAND3X1 NAND3X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_12596_), .B(_12754_), .C(_12749_), .Y(_12755_) );
	AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_12591_), .B(_12595_), .Y(_12756_) );
	OAI21X1 OAI21X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_12752_), .B(_12753_), .C(_12598_), .Y(_12757_) );
	NAND3X1 NAND3X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_12741_), .B(_12748_), .C(_12751_), .Y(_12759_) );
	NAND3X1 NAND3X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_12756_), .B(_12757_), .C(_12759_), .Y(_12760_) );
	NAND3X1 NAND3X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_12760_), .B(_12755_), .C(_12564_), .Y(_12761_) );
	NOR3X1 NOR3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_12517_), .B(_12516_), .C(_12515_), .Y(_12762_) );
	AOI21X1 AOI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_12360_), .B(_12519_), .C(_12762_), .Y(_12763_) );
	AOI21X1 AOI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_12759_), .B(_12757_), .C(_12756_), .Y(_12764_) );
	AOI21X1 AOI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_12749_), .B(_12754_), .C(_12596_), .Y(_12765_) );
	OAI21X1 OAI21X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_12765_), .B(_12764_), .C(_12763_), .Y(_12766_) );
	NAND3X1 NAND3X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_12562_), .B(_12761_), .C(_12766_), .Y(_12767_) );
	OAI21X1 OAI21X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_12765_), .B(_12764_), .C(_12564_), .Y(_12768_) );
	NAND3X1 NAND3X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_12755_), .B(_12760_), .C(_12763_), .Y(_12770_) );
	NAND3X1 NAND3X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12768_), .C(_12770_), .Y(_12771_) );
	NAND3X1 NAND3X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_12767_), .B(_12560_), .C(_12771_), .Y(_12772_) );
	INVX1 INVX1_1809 ( .gnd(gnd), .vdd(vdd), .A(_12560_), .Y(_12773_) );
	AOI21X1 AOI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_12770_), .B(_12768_), .C(_12358_), .Y(_12774_) );
	AOI21X1 AOI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_12766_), .B(_12761_), .C(_12562_), .Y(_12775_) );
	OAI21X1 OAI21X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_12775_), .B(_12774_), .C(_12773_), .Y(_12776_) );
	NAND3X1 NAND3X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .B(_12776_), .C(_12558_), .Y(_12777_) );
	OAI21X1 OAI21X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_12775_), .B(_12774_), .C(_12560_), .Y(_12778_) );
	NAND3X1 NAND3X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_12767_), .B(_12771_), .C(_12773_), .Y(_12779_) );
	NAND3X1 NAND3X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_12536_), .B(_12778_), .C(_12779_), .Y(_12781_) );
	NAND3X1 NAND3X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_12543_), .B(_12781_), .C(_12777_), .Y(_12782_) );
	AOI21X1 AOI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_12546_), .B(_12545_), .C(_12544_), .Y(_12783_) );
	NAND3X1 NAND3X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_12536_), .B(_12772_), .C(_12776_), .Y(_12784_) );
	NAND3X1 NAND3X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_12778_), .B(_12779_), .C(_12558_), .Y(_12785_) );
	NAND3X1 NAND3X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_12784_), .B(_12783_), .C(_12785_), .Y(_12786_) );
	NAND2X1 NAND2X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_12782_), .B(_12786_), .Y(_12787_) );
	XNOR2X1 XNOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_12557_), .B(_12787_), .Y(mulOut_17_) );
	NAND2X1 NAND2X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_12781_), .B(_12777_), .Y(_12788_) );
	NAND3X1 NAND3X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_12543_), .B(_12784_), .C(_12785_), .Y(_12789_) );
	NAND2X1 NAND2X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_12556_), .B(_12789_), .Y(_12791_) );
	OAI21X1 OAI21X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_12543_), .B(_12788_), .C(_12791_), .Y(_12792_) );
	AOI22X1 AOI22X1_287 ( .gnd(gnd), .vdd(vdd), .A(_12548_), .B(_12553_), .C(_12782_), .D(_12786_), .Y(_12793_) );
	AOI21X1 AOI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_12555_), .B(_12793_), .C(_12792_), .Y(_12794_) );
	INVX1 INVX1_1810 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .Y(_12795_) );
	AOI21X1 AOI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_12755_), .B(_12760_), .C(_12564_), .Y(_12796_) );
	OAI21X1 OAI21X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_12358_), .B(_12796_), .C(_12761_), .Y(_12797_) );
	INVX1 INVX1_1811 ( .gnd(gnd), .vdd(vdd), .A(_12587_), .Y(_12798_) );
	AOI21X1 AOI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_12355_), .B(_12590_), .C(_12798_), .Y(_12799_) );
	INVX1 INVX1_1812 ( .gnd(gnd), .vdd(vdd), .A(_12799_), .Y(_12800_) );
	AOI21X1 AOI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_12741_), .B(_12748_), .C(_12598_), .Y(_12802_) );
	OAI21X1 OAI21X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_12756_), .B(_12802_), .C(_12749_), .Y(_12803_) );
	NOR2X1 NOR2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_12347_), .B(_12584_), .Y(_12804_) );
	INVX1 INVX1_1813 ( .gnd(gnd), .vdd(vdd), .A(_12804_), .Y(_12805_) );
	NAND2X1 NAND2X1_2649 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf0), .B(adder_bOperand_18_bF_buf3), .Y(_12806_) );
	INVX1 INVX1_1814 ( .gnd(gnd), .vdd(vdd), .A(_12806_), .Y(_12807_) );
	OAI21X1 OAI21X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_12343_), .B(_12574_), .C(_12573_), .Y(_12808_) );
	NOR2X1 NOR2X1_884 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_12566_), .Y(_12809_) );
	INVX1 INVX1_1815 ( .gnd(gnd), .vdd(vdd), .A(_12809_), .Y(_12810_) );
	NAND2X1 NAND2X1_2650 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .B(adder_bOperand_16_bF_buf1), .Y(_12811_) );
	OAI21X1 OAI21X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_12131_), .C(_12574_), .Y(_12813_) );
	OAI21X1 OAI21X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_12568_), .B(_12811_), .C(_12813_), .Y(_12814_) );
	OR2X2 OR2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_12814_), .B(_12810_), .Y(_12815_) );
	OAI21X1 OAI21X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_12566_), .C(_12814_), .Y(_12816_) );
	NAND2X1 NAND2X1_2651 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf2), .B(adder_bOperand_12_bF_buf2), .Y(_12817_) );
	NOR2X1 NOR2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_12367_), .B(_12817_), .Y(_12818_) );
	AOI21X1 AOI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_12603_), .B(_12601_), .C(_12818_), .Y(_12819_) );
	INVX1 INVX1_1816 ( .gnd(gnd), .vdd(vdd), .A(_12819_), .Y(_12820_) );
	NAND3X1 NAND3X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_12816_), .B(_12820_), .C(_12815_), .Y(_12821_) );
	NOR2X1 NOR2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_12810_), .B(_12814_), .Y(_12822_) );
	AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(adder_bOperand_16_bF_buf0), .Y(_12823_) );
	NAND2X1 NAND2X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_12823_), .B(_12569_), .Y(_12824_) );
	AOI21X1 AOI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_12824_), .B(_12813_), .C(_12809_), .Y(_12825_) );
	OAI21X1 OAI21X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_12825_), .B(_12822_), .C(_12819_), .Y(_12826_) );
	NAND3X1 NAND3X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_12808_), .B(_12826_), .C(_12821_), .Y(_12827_) );
	INVX1 INVX1_1817 ( .gnd(gnd), .vdd(vdd), .A(_12808_), .Y(_12828_) );
	NOR3X1 NOR3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_12819_), .B(_12825_), .C(_12822_), .Y(_12829_) );
	AOI21X1 AOI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_12815_), .B(_12816_), .C(_12820_), .Y(_12830_) );
	OAI21X1 OAI21X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_12829_), .B(_12830_), .C(_12828_), .Y(_12831_) );
	AOI21X1 AOI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_12340_), .C(_12582_), .Y(_12832_) );
	NAND3X1 NAND3X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_12832_), .B(_12827_), .C(_12831_), .Y(_12834_) );
	NAND3X1 NAND3X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_12816_), .B(_12819_), .C(_12815_), .Y(_12835_) );
	OAI21X1 OAI21X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_12825_), .B(_12822_), .C(_12820_), .Y(_12836_) );
	AOI21X1 AOI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_12835_), .B(_12836_), .C(_12828_), .Y(_12837_) );
	AOI21X1 AOI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_12821_), .B(_12826_), .C(_12808_), .Y(_12838_) );
	NAND2X1 NAND2X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_12340_), .B(_12581_), .Y(_12839_) );
	NAND2X1 NAND2X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_12583_), .B(_12839_), .Y(_12840_) );
	OAI21X1 OAI21X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_12837_), .B(_12838_), .C(_12840_), .Y(_12841_) );
	NAND3X1 NAND3X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_12807_), .B(_12834_), .C(_12841_), .Y(_12842_) );
	OAI21X1 OAI21X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_12837_), .B(_12838_), .C(_12832_), .Y(_12843_) );
	NAND3X1 NAND3X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_12827_), .B(_12840_), .C(_12831_), .Y(_12846_) );
	NAND3X1 NAND3X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_12806_), .B(_12843_), .C(_12846_), .Y(_12847_) );
	OAI21X1 OAI21X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_12632_), .B(_12640_), .C(_12642_), .Y(_12848_) );
	NAND3X1 NAND3X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_12842_), .B(_12847_), .C(_12848_), .Y(_12849_) );
	AOI21X1 AOI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_12846_), .B(_12843_), .C(_12806_), .Y(_12850_) );
	AOI21X1 AOI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_12841_), .B(_12834_), .C(_12807_), .Y(_12851_) );
	AOI21X1 AOI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_12599_), .B(_12641_), .C(_12638_), .Y(_12852_) );
	OAI21X1 OAI21X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_12851_), .B(_12850_), .C(_12852_), .Y(_12853_) );
	NAND3X1 NAND3X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_12805_), .B(_12849_), .C(_12853_), .Y(_12854_) );
	NAND3X1 NAND3X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_12842_), .B(_12847_), .C(_12852_), .Y(_12855_) );
	OAI21X1 OAI21X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_12851_), .B(_12850_), .C(_12848_), .Y(_12856_) );
	NAND3X1 NAND3X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_12804_), .B(_12855_), .C(_12856_), .Y(_12857_) );
	NAND2X1 NAND2X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_12857_), .B(_12854_), .Y(_12858_) );
	AOI21X1 AOI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_12734_), .B(_12728_), .C(_12645_), .Y(_12859_) );
	OAI21X1 OAI21X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_12859_), .B(_12744_), .C(_12735_), .Y(_12860_) );
	NAND2X1 NAND2X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_12619_), .B(_12624_), .Y(_12861_) );
	NAND2X1 NAND2X1_2657 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf4), .B(adder_bOperand_14_bF_buf3), .Y(_12862_) );
	INVX1 INVX1_1818 ( .gnd(gnd), .vdd(vdd), .A(_12862_), .Y(_12863_) );
	NAND2X1 NAND2X1_2658 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf4), .B(adder_bOperand_13_bF_buf3), .Y(_12864_) );
	OAI21X1 OAI21X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf1), .B(_17157_), .C(_12602_), .Y(_12865_) );
	OAI21X1 OAI21X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_12817_), .B(_12864_), .C(_12865_), .Y(_12868_) );
	XNOR2X1 XNOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_12868_), .B(_12863_), .Y(_12869_) );
	INVX1 INVX1_1819 ( .gnd(gnd), .vdd(vdd), .A(_12376_), .Y(_12870_) );
	AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf1), .B(adder_bOperand_10_bF_buf1), .Y(_12871_) );
	AOI22X1 AOI22X1_288 ( .gnd(gnd), .vdd(vdd), .A(_12870_), .B(_12871_), .C(_12608_), .D(_12612_), .Y(_12872_) );
	INVX1 INVX1_1820 ( .gnd(gnd), .vdd(vdd), .A(_12872_), .Y(_12873_) );
	NAND2X1 NAND2X1_2659 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf3), .B(adder_bOperand_11_bF_buf3), .Y(_12874_) );
	INVX1 INVX1_1821 ( .gnd(gnd), .vdd(vdd), .A(_12874_), .Y(_12875_) );
	AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf2), .B(adder_bOperand_10_bF_buf0), .Y(_12876_) );
	NAND2X1 NAND2X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_12610_), .B(_12876_), .Y(_12877_) );
	NAND2X1 NAND2X1_2661 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf0), .B(adder_bOperand_10_bF_buf4), .Y(_12879_) );
	OAI21X1 OAI21X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf2), .B(_17025__bF_buf3), .C(_12879_), .Y(_12880_) );
	NAND3X1 NAND3X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_12875_), .B(_12880_), .C(_12877_), .Y(_12881_) );
	NAND2X1 NAND2X1_2662 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf1), .B(adder_bOperand_9_bF_buf2), .Y(_12882_) );
	NOR2X1 NOR2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_12879_), .B(_12882_), .Y(_12883_) );
	AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_12879_), .B(_12882_), .Y(_12884_) );
	OAI21X1 OAI21X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_12883_), .B(_12884_), .C(_12874_), .Y(_12885_) );
	NAND3X1 NAND3X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_12885_), .C(_12873_), .Y(_12886_) );
	NOR3X1 NOR3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_12874_), .B(_12883_), .C(_12884_), .Y(_12887_) );
	AOI21X1 AOI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_12877_), .B(_12880_), .C(_12875_), .Y(_12888_) );
	OAI21X1 OAI21X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_12888_), .B(_12887_), .C(_12872_), .Y(_12890_) );
	NAND3X1 NAND3X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_12869_), .B(_12890_), .C(_12886_), .Y(_12891_) );
	XNOR2X1 XNOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_12868_), .B(_12862_), .Y(_12892_) );
	OAI21X1 OAI21X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_12888_), .B(_12887_), .C(_12873_), .Y(_12893_) );
	NAND3X1 NAND3X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_12881_), .B(_12872_), .C(_12885_), .Y(_12894_) );
	NAND3X1 NAND3X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_12894_), .B(_12892_), .C(_12893_), .Y(_12895_) );
	AOI21X1 AOI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_12653_), .B(_12658_), .C(_12663_), .Y(_12896_) );
	OAI21X1 OAI21X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_12646_), .B(_12896_), .C(_12664_), .Y(_12897_) );
	AOI21X1 AOI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_12891_), .B(_12895_), .C(_12897_), .Y(_12898_) );
	AOI21X1 AOI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_12893_), .B(_12894_), .C(_12892_), .Y(_12899_) );
	AOI21X1 AOI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_12886_), .B(_12890_), .C(_12869_), .Y(_12901_) );
	NOR3X1 NOR3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .B(_12665_), .C(_12666_), .Y(_12902_) );
	AOI21X1 AOI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_12667_), .B(_12669_), .C(_12902_), .Y(_12903_) );
	NOR3X1 NOR3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(_12901_), .C(_12903_), .Y(_12904_) );
	OAI21X1 OAI21X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .B(_12904_), .C(_12861_), .Y(_12905_) );
	INVX1 INVX1_1822 ( .gnd(gnd), .vdd(vdd), .A(_12861_), .Y(_12906_) );
	INVX1 INVX1_1823 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .Y(_12907_) );
	NAND3X1 NAND3X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_12891_), .B(_12895_), .C(_12897_), .Y(_12908_) );
	NAND3X1 NAND3X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_12906_), .B(_12908_), .C(_12907_), .Y(_12909_) );
	NAND2X1 NAND2X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_12909_), .B(_12905_), .Y(_12910_) );
	AOI21X1 AOI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_12713_), .B(_12720_), .C(_12676_), .Y(_12912_) );
	OAI21X1 OAI21X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_12731_), .B(_12912_), .C(_12721_), .Y(_12913_) );
	NAND2X1 NAND2X1_2664 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf0), .B(aOperand_frameOut_11_bF_buf3), .Y(_12914_) );
	OAI21X1 OAI21X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_12416_), .B(_12914_), .C(_12653_), .Y(_12915_) );
	NAND2X1 NAND2X1_2665 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf3), .B(aOperand_frameOut_10_bF_buf0), .Y(_12916_) );
	INVX1 INVX1_1824 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .Y(_12917_) );
	AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf0), .B(aOperand_frameOut_12_bF_buf3), .Y(_12918_) );
	NAND2X1 NAND2X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_12649_), .B(_12918_), .Y(_12919_) );
	OAI21X1 OAI21X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf1), .B(_17236__bF_buf2), .C(_12914_), .Y(_12920_) );
	NAND3X1 NAND3X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_12917_), .B(_12920_), .C(_12919_), .Y(_12921_) );
	NAND3X1 NAND3X1_2751 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(aOperand_frameOut_12_bF_buf2), .C(_12914_), .Y(_12923_) );
	NAND2X1 NAND2X1_2667 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf4), .B(aOperand_frameOut_12_bF_buf1), .Y(_12924_) );
	NAND3X1 NAND3X1_2752 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(aOperand_frameOut_11_bF_buf2), .C(_12924_), .Y(_12925_) );
	NAND3X1 NAND3X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_12916_), .B(_12923_), .C(_12925_), .Y(_12926_) );
	OAI21X1 OAI21X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_12677_), .B(_12688_), .C(_12680_), .Y(_12927_) );
	AOI21X1 AOI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_12921_), .B(_12926_), .C(_12927_), .Y(_12928_) );
	AOI21X1 AOI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_12923_), .B(_12925_), .C(_12916_), .Y(_12929_) );
	AOI21X1 AOI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_12919_), .B(_12920_), .C(_12917_), .Y(_12930_) );
	AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf5), .B(aOperand_frameOut_14_bF_buf4), .Y(_12931_) );
	AOI22X1 AOI22X1_289 ( .gnd(gnd), .vdd(vdd), .A(_12446_), .B(_12931_), .C(_12685_), .D(_12683_), .Y(_12932_) );
	NOR3X1 NOR3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_12932_), .B(_12929_), .C(_12930_), .Y(_12934_) );
	OAI21X1 OAI21X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12934_), .C(_12915_), .Y(_12935_) );
	AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_12653_), .B(_12650_), .Y(_12936_) );
	OAI21X1 OAI21X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_12929_), .B(_12930_), .C(_12932_), .Y(_12937_) );
	NAND3X1 NAND3X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_12921_), .B(_12926_), .C(_12927_), .Y(_12938_) );
	NAND3X1 NAND3X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_12937_), .B(_12938_), .C(_12936_), .Y(_12939_) );
	NAND2X1 NAND2X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_12939_), .B(_12935_), .Y(_12940_) );
	AOI21X1 AOI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_12704_), .B(_12700_), .C(_12691_), .Y(_12941_) );
	OAI21X1 OAI21X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_12717_), .B(_12941_), .C(_12705_), .Y(_12942_) );
	NAND2X1 NAND2X1_2669 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf2), .B(aOperand_frameOut_13_bF_buf1), .Y(_12943_) );
	AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf0), .B(aOperand_frameOut_15_bF_buf1), .Y(_12945_) );
	NAND2X1 NAND2X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_12931_), .B(_12945_), .Y(_12946_) );
	NAND2X1 NAND2X1_2671 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf5), .B(aOperand_frameOut_15_bF_buf0), .Y(_12947_) );
	NAND2X1 NAND2X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_12686_), .B(_12947_), .Y(_12948_) );
	NAND3X1 NAND3X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(_12948_), .C(_12946_), .Y(_12949_) );
	INVX1 INVX1_1825 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .Y(_12950_) );
	OAI21X1 OAI21X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_12039_), .C(_12945_), .Y(_12951_) );
	OAI21X1 OAI21X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf1), .B(_12233_), .C(_12931_), .Y(_12952_) );
	NAND3X1 NAND3X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_12951_), .C(_12952_), .Y(_12953_) );
	NAND2X1 NAND2X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_12949_), .B(_12953_), .Y(_12954_) );
	OAI21X1 OAI21X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_12693_), .B(_12702_), .C(_12697_), .Y(_12956_) );
	NAND2X1 NAND2X1_2674 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf0), .B(aOperand_frameOut_16_bF_buf0), .Y(_12957_) );
	INVX1 INVX1_1826 ( .gnd(gnd), .vdd(vdd), .A(_12957_), .Y(_12958_) );
	AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf0), .B(aOperand_frameOut_18_bF_buf0), .Y(_12959_) );
	NAND2X1 NAND2X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_12696_), .B(_12959_), .Y(_12960_) );
	NAND2X1 NAND2X1_2676 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf6), .B(aOperand_frameOut_17_bF_buf3), .Y(_12961_) );
	NAND2X1 NAND2X1_2677 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_18_bF_buf4), .Y(_12962_) );
	NAND2X1 NAND2X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_12961_), .B(_12962_), .Y(_12963_) );
	NAND3X1 NAND3X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_12958_), .B(_12963_), .C(_12960_), .Y(_12964_) );
	NAND3X1 NAND3X1_2759 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_18_bF_buf3), .C(_12961_), .Y(_12965_) );
	NAND3X1 NAND3X1_2760 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(aOperand_frameOut_17_bF_buf2), .C(_12962_), .Y(_12967_) );
	NAND3X1 NAND3X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_12957_), .B(_12965_), .C(_12967_), .Y(_12968_) );
	NAND3X1 NAND3X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_12964_), .B(_12968_), .C(_12956_), .Y(_12969_) );
	AOI21X1 AOI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_12694_), .B(_12699_), .C(_12701_), .Y(_12970_) );
	AOI21X1 AOI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_12965_), .B(_12967_), .C(_12957_), .Y(_12971_) );
	AOI21X1 AOI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_12960_), .B(_12963_), .C(_12958_), .Y(_12972_) );
	OAI21X1 OAI21X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_12971_), .B(_12972_), .C(_12970_), .Y(_12973_) );
	NAND3X1 NAND3X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_12954_), .B(_12969_), .C(_12973_), .Y(_12974_) );
	NAND3X1 NAND3X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_12950_), .B(_12948_), .C(_12946_), .Y(_12975_) );
	NAND3X1 NAND3X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(_12951_), .C(_12952_), .Y(_12976_) );
	NAND2X1 NAND2X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_12975_), .B(_12976_), .Y(_12978_) );
	OAI21X1 OAI21X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_12971_), .B(_12972_), .C(_12956_), .Y(_12979_) );
	NAND3X1 NAND3X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_12968_), .B(_12970_), .C(_12964_), .Y(_12980_) );
	NAND3X1 NAND3X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_12978_), .B(_12980_), .C(_12979_), .Y(_12981_) );
	NAND3X1 NAND3X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_12981_), .C(_12942_), .Y(_12982_) );
	NOR3X1 NOR3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_12706_), .B(_12711_), .C(_12710_), .Y(_12983_) );
	AOI21X1 AOI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_12690_), .B(_12712_), .C(_12983_), .Y(_12984_) );
	AOI21X1 AOI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_12979_), .B(_12980_), .C(_12978_), .Y(_12985_) );
	AOI21X1 AOI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_12973_), .B(_12969_), .C(_12954_), .Y(_12986_) );
	OAI21X1 OAI21X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_12985_), .B(_12986_), .C(_12984_), .Y(_12987_) );
	NAND3X1 NAND3X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_12982_), .B(_12940_), .C(_12987_), .Y(_12989_) );
	NAND3X1 NAND3X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(_12937_), .C(_12938_), .Y(_12990_) );
	OAI21X1 OAI21X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12934_), .C(_12936_), .Y(_12991_) );
	NAND2X1 NAND2X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_12990_), .B(_12991_), .Y(_12992_) );
	OAI21X1 OAI21X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_12985_), .B(_12986_), .C(_12942_), .Y(_12993_) );
	NAND3X1 NAND3X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_12981_), .C(_12984_), .Y(_12994_) );
	NAND3X1 NAND3X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_12992_), .B(_12994_), .C(_12993_), .Y(_12995_) );
	NAND3X1 NAND3X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_12989_), .B(_12995_), .C(_12913_), .Y(_12996_) );
	NAND2X1 NAND2X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_12713_), .B(_12720_), .Y(_12997_) );
	NOR2X1 NOR2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_12723_), .B(_12997_), .Y(_12998_) );
	AOI21X1 AOI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_12674_), .B(_12727_), .C(_12998_), .Y(_13000_) );
	AOI21X1 AOI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_12993_), .B(_12994_), .C(_12992_), .Y(_13001_) );
	AOI21X1 AOI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_12987_), .B(_12982_), .C(_12940_), .Y(_13002_) );
	OAI21X1 OAI21X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_13001_), .B(_13002_), .C(_13000_), .Y(_13003_) );
	NAND3X1 NAND3X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_12996_), .B(_13003_), .C(_12910_), .Y(_13004_) );
	NAND3X1 NAND3X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_12861_), .B(_12908_), .C(_12907_), .Y(_13005_) );
	OAI21X1 OAI21X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .B(_12904_), .C(_12906_), .Y(_13006_) );
	NAND2X1 NAND2X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_13005_), .B(_13006_), .Y(_13007_) );
	OAI21X1 OAI21X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_13001_), .B(_13002_), .C(_12913_), .Y(_13008_) );
	NAND3X1 NAND3X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_12989_), .B(_12995_), .C(_13000_), .Y(_13009_) );
	NAND3X1 NAND3X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_13008_), .B(_13009_), .C(_13007_), .Y(_13011_) );
	NAND3X1 NAND3X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_13004_), .B(_13011_), .C(_12860_), .Y(_13012_) );
	INVX1 INVX1_1827 ( .gnd(gnd), .vdd(vdd), .A(_12735_), .Y(_13013_) );
	AOI21X1 AOI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_12644_), .B(_12740_), .C(_13013_), .Y(_13014_) );
	AOI21X1 AOI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_13009_), .B(_13008_), .C(_13007_), .Y(_13015_) );
	AOI22X1 AOI22X1_290 ( .gnd(gnd), .vdd(vdd), .A(_13005_), .B(_13006_), .C(_12996_), .D(_13003_), .Y(_13016_) );
	OAI21X1 OAI21X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_13016_), .B(_13015_), .C(_13014_), .Y(_13017_) );
	NAND3X1 NAND3X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_13012_), .B(_13017_), .C(_12858_), .Y(_13018_) );
	NAND3X1 NAND3X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_12804_), .B(_12849_), .C(_12853_), .Y(_13019_) );
	NAND3X1 NAND3X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_12805_), .B(_12855_), .C(_12856_), .Y(_13020_) );
	NAND2X1 NAND2X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_13020_), .B(_13019_), .Y(_13022_) );
	OAI21X1 OAI21X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_13016_), .B(_13015_), .C(_12860_), .Y(_13023_) );
	NAND3X1 NAND3X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_13004_), .B(_13011_), .C(_13014_), .Y(_13024_) );
	NAND3X1 NAND3X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_13023_), .B(_13024_), .C(_13022_), .Y(_13025_) );
	NAND3X1 NAND3X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_13018_), .B(_13025_), .C(_12803_), .Y(_13026_) );
	NOR3X1 NOR3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_12752_), .B(_12753_), .C(_12751_), .Y(_13027_) );
	AOI21X1 AOI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_12596_), .B(_12754_), .C(_13027_), .Y(_13028_) );
	AOI21X1 AOI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_13024_), .B(_13023_), .C(_13022_), .Y(_13029_) );
	AOI21X1 AOI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_13017_), .B(_13012_), .C(_12858_), .Y(_13030_) );
	OAI21X1 OAI21X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_13029_), .B(_13030_), .C(_13028_), .Y(_13031_) );
	NAND3X1 NAND3X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_12800_), .B(_13026_), .C(_13031_), .Y(_13033_) );
	OAI21X1 OAI21X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_13030_), .B(_13029_), .C(_12803_), .Y(_13034_) );
	NAND3X1 NAND3X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_13018_), .B(_13025_), .C(_13028_), .Y(_13035_) );
	NAND3X1 NAND3X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_12799_), .B(_13034_), .C(_13035_), .Y(_13036_) );
	NAND3X1 NAND3X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_13033_), .B(_13036_), .C(_12797_), .Y(_13037_) );
	INVX1 INVX1_1828 ( .gnd(gnd), .vdd(vdd), .A(_12761_), .Y(_13038_) );
	AOI21X1 AOI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_12562_), .B(_12766_), .C(_13038_), .Y(_13039_) );
	AOI21X1 AOI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_13035_), .B(_13034_), .C(_12799_), .Y(_13040_) );
	AOI21X1 AOI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_13031_), .B(_13026_), .C(_12800_), .Y(_13041_) );
	OAI21X1 OAI21X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_13041_), .B(_13040_), .C(_13039_), .Y(_13042_) );
	NAND3X1 NAND3X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_13037_), .B(_13042_), .C(_12795_), .Y(_13044_) );
	OAI21X1 OAI21X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_13041_), .B(_13040_), .C(_12797_), .Y(_13045_) );
	NAND3X1 NAND3X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_13033_), .B(_13036_), .C(_13039_), .Y(_13046_) );
	NAND3X1 NAND3X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .B(_13045_), .C(_13046_), .Y(_13047_) );
	NAND3X1 NAND3X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_13047_), .B(_13044_), .C(_12777_), .Y(_13048_) );
	AOI21X1 AOI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_12779_), .B(_12778_), .C(_12536_), .Y(_13049_) );
	NAND3X1 NAND3X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .B(_13037_), .C(_13042_), .Y(_13050_) );
	NAND3X1 NAND3X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_13045_), .B(_13046_), .C(_12795_), .Y(_13051_) );
	NAND3X1 NAND3X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_13050_), .B(_13051_), .C(_13049_), .Y(_13052_) );
	NAND2X1 NAND2X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_13048_), .B(_13052_), .Y(_13053_) );
	XNOR2X1 XNOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_12794_), .B(_13053_), .Y(mulOut_18_) );
	NAND3X1 NAND3X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_13047_), .B(_13044_), .C(_13049_), .Y(_13055_) );
	INVX1 INVX1_1829 ( .gnd(gnd), .vdd(vdd), .A(_13053_), .Y(_13056_) );
	OAI21X1 OAI21X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_13056_), .B(_12794_), .C(_13055_), .Y(_13057_) );
	AOI21X1 AOI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_13046_), .B(_13045_), .C(_12772_), .Y(_13058_) );
	AOI21X1 AOI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_13018_), .B(_13025_), .C(_12803_), .Y(_13059_) );
	OAI21X1 OAI21X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_12799_), .B(_13059_), .C(_13026_), .Y(_13060_) );
	NAND2X1 NAND2X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_12849_), .B(_13019_), .Y(_13061_) );
	INVX1 INVX1_1830 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .Y(_13062_) );
	AOI21X1 AOI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_13004_), .B(_13011_), .C(_12860_), .Y(_13063_) );
	OAI21X1 OAI21X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_13063_), .B(_13022_), .C(_13012_), .Y(_13064_) );
	NAND2X1 NAND2X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_12834_), .B(_12842_), .Y(_13065_) );
	NAND2X1 NAND2X1_2687 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf4), .B(adder_bOperand_19_bF_buf2), .Y(_13066_) );
	INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_19_bF_buf1), .Y(_13067_) );
	NAND2X1 NAND2X1_2688 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf3), .B(adder_bOperand_18_bF_buf2), .Y(_13068_) );
	OAI21X1 OAI21X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf1), .B(_13067_), .C(_13068_), .Y(_13069_) );
	OAI21X1 OAI21X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_12806_), .B(_13066_), .C(_13069_), .Y(_13070_) );
	INVX1 INVX1_1831 ( .gnd(gnd), .vdd(vdd), .A(_13070_), .Y(_13071_) );
	OAI21X1 OAI21X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_12828_), .B(_12830_), .C(_12821_), .Y(_13072_) );
	OAI21X1 OAI21X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_12810_), .B(_12814_), .C(_12824_), .Y(_13073_) );
	NAND2X1 NAND2X1_2689 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf2), .B(adder_bOperand_17_bF_buf3), .Y(_13075_) );
	INVX1 INVX1_1832 ( .gnd(gnd), .vdd(vdd), .A(_13075_), .Y(_13076_) );
	AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .B(adder_bOperand_15_bF_buf2), .Y(_13077_) );
	NAND2X1 NAND2X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_12823_), .B(_13077_), .Y(_13078_) );
	OAI21X1 OAI21X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf1), .B(_12131_), .C(_12811_), .Y(_13079_) );
	NAND3X1 NAND3X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_13076_), .B(_13079_), .C(_13078_), .Y(_13080_) );
	OAI21X1 OAI21X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_12342_), .C(_13077_), .Y(_13081_) );
	OAI21X1 OAI21X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf0), .B(_12131_), .C(_12823_), .Y(_13082_) );
	NAND3X1 NAND3X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_13075_), .B(_13081_), .C(_13082_), .Y(_13083_) );
	NAND2X1 NAND2X1_2691 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf3), .B(adder_bOperand_12_bF_buf1), .Y(_13084_) );
	AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_12602_), .B(_13084_), .Y(_13086_) );
	OAI22X1 OAI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(_12817_), .B(_12864_), .C(_12862_), .D(_13086_), .Y(_13087_) );
	NAND3X1 NAND3X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_13080_), .B(_13083_), .C(_13087_), .Y(_13088_) );
	AOI21X1 AOI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_13081_), .B(_13082_), .C(_13075_), .Y(_13089_) );
	AOI21X1 AOI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_13078_), .B(_13079_), .C(_13076_), .Y(_13090_) );
	NOR2X1 NOR2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_12602_), .B(_13084_), .Y(_13091_) );
	AOI21X1 AOI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_12865_), .B(_12863_), .C(_13091_), .Y(_13092_) );
	OAI21X1 OAI21X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_13090_), .B(_13089_), .C(_13092_), .Y(_13093_) );
	NAND3X1 NAND3X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_13073_), .B(_13088_), .C(_13093_), .Y(_13094_) );
	AOI21X1 AOI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_13093_), .B(_13088_), .C(_13073_), .Y(_13095_) );
	INVX1 INVX1_1833 ( .gnd(gnd), .vdd(vdd), .A(_13095_), .Y(_13097_) );
	NAND3X1 NAND3X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_13094_), .B(_13097_), .C(_13072_), .Y(_13098_) );
	AOI21X1 AOI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_12826_), .B(_12808_), .C(_12829_), .Y(_13099_) );
	INVX1 INVX1_1834 ( .gnd(gnd), .vdd(vdd), .A(_13094_), .Y(_13100_) );
	OAI21X1 OAI21X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_13095_), .B(_13100_), .C(_13099_), .Y(_13101_) );
	NAND3X1 NAND3X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_13071_), .B(_13101_), .C(_13098_), .Y(_13102_) );
	OAI21X1 OAI21X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_13095_), .B(_13100_), .C(_13072_), .Y(_13103_) );
	NAND3X1 NAND3X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_13099_), .B(_13094_), .C(_13097_), .Y(_13104_) );
	NAND3X1 NAND3X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_13070_), .B(_13104_), .C(_13103_), .Y(_13105_) );
	OAI21X1 OAI21X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_12898_), .B(_12906_), .C(_12908_), .Y(_13106_) );
	NAND3X1 NAND3X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_13106_), .B(_13105_), .C(_13102_), .Y(_13108_) );
	AOI21X1 AOI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_13103_), .B(_13104_), .C(_13070_), .Y(_13109_) );
	AOI21X1 AOI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_13098_), .B(_13101_), .C(_13071_), .Y(_13110_) );
	AOI21X1 AOI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_12907_), .B(_12861_), .C(_12904_), .Y(_13111_) );
	OAI21X1 OAI21X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_13109_), .B(_13110_), .C(_13111_), .Y(_13112_) );
	NAND3X1 NAND3X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_13065_), .B(_13108_), .C(_13112_), .Y(_13113_) );
	AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_12842_), .B(_12834_), .Y(_13114_) );
	NAND3X1 NAND3X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_13105_), .B(_13102_), .C(_13111_), .Y(_13115_) );
	OAI21X1 OAI21X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_13109_), .B(_13110_), .C(_13106_), .Y(_13116_) );
	NAND3X1 NAND3X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_13114_), .B(_13116_), .C(_13115_), .Y(_13117_) );
	NAND2X1 NAND2X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_13113_), .B(_13117_), .Y(_13119_) );
	AOI21X1 AOI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_12995_), .B(_12989_), .C(_12913_), .Y(_13120_) );
	OAI21X1 OAI21X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_13120_), .B(_13007_), .C(_12996_), .Y(_13121_) );
	NAND2X1 NAND2X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_12886_), .B(_12891_), .Y(_13122_) );
	NAND2X1 NAND2X1_2694 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf1), .B(adder_bOperand_14_bF_buf2), .Y(_13123_) );
	NAND2X1 NAND2X1_2695 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf2), .B(adder_bOperand_13_bF_buf2), .Y(_13124_) );
	OAI21X1 OAI21X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_17157_), .C(_12864_), .Y(_13125_) );
	OAI21X1 OAI21X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_13084_), .B(_13124_), .C(_13125_), .Y(_13126_) );
	XNOR2X1 XNOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_13126_), .B(_13123_), .Y(_13127_) );
	OAI21X1 OAI21X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_12874_), .B(_12884_), .C(_12877_), .Y(_13128_) );
	NAND2X1 NAND2X1_2696 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf4), .B(adder_bOperand_11_bF_buf2), .Y(_13130_) );
	AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf4), .B(adder_bOperand_9_bF_buf1), .Y(_13131_) );
	OAI21X1 OAI21X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf1), .B(_16887_), .C(_13131_), .Y(_13132_) );
	OAI21X1 OAI21X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_17025__bF_buf2), .C(_12876_), .Y(_13133_) );
	AOI21X1 AOI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_13132_), .B(_13133_), .C(_13130_), .Y(_13134_) );
	INVX1 INVX1_1835 ( .gnd(gnd), .vdd(vdd), .A(_13130_), .Y(_13135_) );
	NAND2X1 NAND2X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_12876_), .B(_13131_), .Y(_13136_) );
	NAND2X1 NAND2X1_2698 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf0), .B(adder_bOperand_10_bF_buf3), .Y(_13137_) );
	OAI21X1 OAI21X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_17025__bF_buf1), .C(_13137_), .Y(_13138_) );
	AOI21X1 AOI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_13136_), .B(_13138_), .C(_13135_), .Y(_13139_) );
	OAI21X1 OAI21X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_13139_), .B(_13134_), .C(_13128_), .Y(_13141_) );
	AOI21X1 AOI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_12880_), .B(_12875_), .C(_12883_), .Y(_13142_) );
	NAND3X1 NAND3X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_13135_), .B(_13138_), .C(_13136_), .Y(_13143_) );
	NAND2X1 NAND2X1_2699 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf3), .B(adder_bOperand_9_bF_buf0), .Y(_13144_) );
	NOR2X1 NOR2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_13137_), .B(_13144_), .Y(_13145_) );
	AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_13137_), .B(_13144_), .Y(_13146_) );
	OAI21X1 OAI21X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_13145_), .B(_13146_), .C(_13130_), .Y(_13147_) );
	NAND3X1 NAND3X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_13143_), .B(_13142_), .C(_13147_), .Y(_13148_) );
	AOI21X1 AOI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_13141_), .B(_13148_), .C(_13127_), .Y(_13149_) );
	INVX1 INVX1_1836 ( .gnd(gnd), .vdd(vdd), .A(_13123_), .Y(_13150_) );
	XNOR2X1 XNOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_13126_), .B(_13150_), .Y(_13152_) );
	NAND3X1 NAND3X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_13143_), .B(_13128_), .C(_13147_), .Y(_13153_) );
	OAI21X1 OAI21X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_13139_), .B(_13134_), .C(_13142_), .Y(_13154_) );
	AOI21X1 AOI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_13154_), .B(_13153_), .C(_13152_), .Y(_13155_) );
	AOI21X1 AOI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(_12937_), .C(_12934_), .Y(_13156_) );
	OAI21X1 OAI21X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_13149_), .B(_13155_), .C(_13156_), .Y(_13157_) );
	NAND3X1 NAND3X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_13153_), .B(_13154_), .C(_13152_), .Y(_13158_) );
	NAND3X1 NAND3X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_13148_), .B(_13141_), .C(_13127_), .Y(_13159_) );
	OAI21X1 OAI21X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12936_), .C(_12938_), .Y(_13160_) );
	NAND3X1 NAND3X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_13159_), .B(_13158_), .C(_13160_), .Y(_13161_) );
	NAND3X1 NAND3X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .B(_13161_), .C(_13157_), .Y(_13163_) );
	INVX1 INVX1_1837 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .Y(_13164_) );
	AOI21X1 AOI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_13158_), .B(_13159_), .C(_13160_), .Y(_13165_) );
	NOR3X1 NOR3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_13149_), .B(_13155_), .C(_13156_), .Y(_13166_) );
	OAI21X1 OAI21X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_13165_), .B(_13166_), .C(_13164_), .Y(_13167_) );
	NAND2X1 NAND2X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_13163_), .B(_13167_), .Y(_13168_) );
	AOI21X1 AOI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_12974_), .B(_12981_), .C(_12942_), .Y(_13169_) );
	OAI21X1 OAI21X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_13169_), .B(_12992_), .C(_12982_), .Y(_13170_) );
	NAND2X1 NAND2X1_2701 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf4), .B(aOperand_frameOut_12_bF_buf0), .Y(_13171_) );
	OAI21X1 OAI21X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_12656_), .B(_13171_), .C(_12921_), .Y(_13172_) );
	NAND2X1 NAND2X1_2702 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf2), .B(aOperand_frameOut_11_bF_buf1), .Y(_13174_) );
	NAND3X1 NAND3X1_2816 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf3), .B(aOperand_frameOut_13_bF_buf0), .C(_13171_), .Y(_13175_) );
	NAND2X1 NAND2X1_2703 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf2), .B(aOperand_frameOut_13_bF_buf4), .Y(_13176_) );
	NAND3X1 NAND3X1_2817 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf3), .B(aOperand_frameOut_12_bF_buf4), .C(_13176_), .Y(_13177_) );
	AOI21X1 AOI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_13175_), .B(_13177_), .C(_13174_), .Y(_13178_) );
	INVX1 INVX1_1838 ( .gnd(gnd), .vdd(vdd), .A(_13174_), .Y(_13179_) );
	AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf2), .B(aOperand_frameOut_13_bF_buf3), .Y(_13180_) );
	NAND2X1 NAND2X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_12918_), .B(_13180_), .Y(_13181_) );
	OAI21X1 OAI21X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf0), .B(_11858_), .C(_13171_), .Y(_13182_) );
	AOI21X1 AOI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_13181_), .B(_13182_), .C(_13179_), .Y(_13183_) );
	AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .B(aOperand_frameOut_15_bF_buf4), .Y(_13185_) );
	AOI22X1 AOI22X1_291 ( .gnd(gnd), .vdd(vdd), .A(_12679_), .B(_13185_), .C(_12950_), .D(_12948_), .Y(_13186_) );
	OAI21X1 OAI21X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_13178_), .B(_13183_), .C(_13186_), .Y(_13187_) );
	NAND3X1 NAND3X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_13179_), .B(_13182_), .C(_13181_), .Y(_13188_) );
	NAND3X1 NAND3X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_13174_), .B(_13175_), .C(_13177_), .Y(_13189_) );
	INVX1 INVX1_1839 ( .gnd(gnd), .vdd(vdd), .A(_13186_), .Y(_13190_) );
	NAND3X1 NAND3X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_13188_), .B(_13189_), .C(_13190_), .Y(_13191_) );
	NAND3X1 NAND3X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_13172_), .B(_13187_), .C(_13191_), .Y(_13192_) );
	AOI21X1 AOI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_12649_), .B(_12918_), .C(_12929_), .Y(_13193_) );
	AOI21X1 AOI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_13188_), .B(_13189_), .C(_13190_), .Y(_13194_) );
	NOR3X1 NOR3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_13186_), .B(_13178_), .C(_13183_), .Y(_13196_) );
	OAI21X1 OAI21X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_13194_), .B(_13196_), .C(_13193_), .Y(_13197_) );
	NAND2X1 NAND2X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_13192_), .B(_13197_), .Y(_13198_) );
	AOI21X1 AOI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_12964_), .B(_12968_), .C(_12956_), .Y(_13199_) );
	OAI21X1 OAI21X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_12978_), .B(_13199_), .C(_12969_), .Y(_13200_) );
	NAND2X1 NAND2X1_2706 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf1), .B(aOperand_frameOut_14_bF_buf3), .Y(_13201_) );
	AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .B(aOperand_frameOut_16_bF_buf4), .Y(_13202_) );
	NAND2X1 NAND2X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_13185_), .B(_13202_), .Y(_13203_) );
	NAND2X1 NAND2X1_2708 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf3), .B(aOperand_frameOut_15_bF_buf3), .Y(_13204_) );
	NAND2X1 NAND2X1_2709 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf3), .B(aOperand_frameOut_16_bF_buf3), .Y(_13205_) );
	NAND2X1 NAND2X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_13204_), .B(_13205_), .Y(_13207_) );
	NAND3X1 NAND3X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_13201_), .B(_13207_), .C(_13203_), .Y(_13208_) );
	INVX1 INVX1_1840 ( .gnd(gnd), .vdd(vdd), .A(_13201_), .Y(_13209_) );
	OAI21X1 OAI21X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_12233_), .C(_13202_), .Y(_13210_) );
	OAI21X1 OAI21X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf0), .B(_12461_), .C(_13185_), .Y(_13211_) );
	NAND3X1 NAND3X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_13209_), .B(_13210_), .C(_13211_), .Y(_13212_) );
	AOI22X1 AOI22X1_292 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_18_bF_buf2), .C(adder_bOperand_1_bF_buf4), .D(aOperand_frameOut_17_bF_buf1), .Y(_13213_) );
	OAI21X1 OAI21X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_12957_), .B(_13213_), .C(_12960_), .Y(_13214_) );
	NAND2X1 NAND2X1_2711 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf5), .B(aOperand_frameOut_17_bF_buf0), .Y(_13215_) );
	NAND2X1 NAND2X1_2712 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf3), .B(aOperand_frameOut_18_bF_buf1), .Y(_13216_) );
	NAND3X1 NAND3X1_2824 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(aOperand_frameOut_19_bF_buf0), .C(_13216_), .Y(_13218_) );
	NAND2X1 NAND2X1_2713 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .B(aOperand_frameOut_19_bF_buf4), .Y(_13219_) );
	NAND3X1 NAND3X1_2825 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .B(aOperand_frameOut_18_bF_buf0), .C(_13219_), .Y(_13220_) );
	AOI21X1 AOI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_13218_), .B(_13220_), .C(_13215_), .Y(_13221_) );
	AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(aOperand_frameOut_19_bF_buf3), .Y(_13222_) );
	NAND2X1 NAND2X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_12959_), .B(_13222_), .Y(_13223_) );
	INVX4 INVX4_20 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_19_bF_buf2), .Y(_13224_) );
	OAI21X1 OAI21X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf3), .B(_13224_), .C(_13216_), .Y(_13225_) );
	AOI22X1 AOI22X1_293 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .B(aOperand_frameOut_17_bF_buf4), .C(_13225_), .D(_13223_), .Y(_13226_) );
	OAI21X1 OAI21X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_13221_), .B(_13226_), .C(_13214_), .Y(_13227_) );
	AOI22X1 AOI22X1_294 ( .gnd(gnd), .vdd(vdd), .A(_12696_), .B(_12959_), .C(_12958_), .D(_12963_), .Y(_13229_) );
	INVX1 INVX1_1841 ( .gnd(gnd), .vdd(vdd), .A(_13215_), .Y(_13230_) );
	NAND3X1 NAND3X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_13230_), .B(_13225_), .C(_13223_), .Y(_13231_) );
	NAND3X1 NAND3X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_13215_), .B(_13218_), .C(_13220_), .Y(_13232_) );
	NAND3X1 NAND3X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_13229_), .B(_13232_), .C(_13231_), .Y(_13233_) );
	AOI22X1 AOI22X1_295 ( .gnd(gnd), .vdd(vdd), .A(_13208_), .B(_13212_), .C(_13233_), .D(_13227_), .Y(_13234_) );
	NAND2X1 NAND2X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_13208_), .B(_13212_), .Y(_13235_) );
	NAND3X1 NAND3X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_13232_), .B(_13214_), .C(_13231_), .Y(_13236_) );
	OAI21X1 OAI21X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_13221_), .B(_13226_), .C(_13229_), .Y(_13237_) );
	AOI21X1 AOI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_13237_), .B(_13236_), .C(_13235_), .Y(_13238_) );
	OAI21X1 OAI21X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_13234_), .B(_13238_), .C(_13200_), .Y(_13240_) );
	NOR3X1 NOR3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_12970_), .B(_12971_), .C(_12972_), .Y(_13241_) );
	AOI21X1 AOI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_12954_), .B(_12973_), .C(_13241_), .Y(_13242_) );
	NAND3X1 NAND3X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_13235_), .B(_13236_), .C(_13237_), .Y(_13243_) );
	NAND3X1 NAND3X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_13209_), .B(_13207_), .C(_13203_), .Y(_13244_) );
	NAND3X1 NAND3X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_13201_), .B(_13210_), .C(_13211_), .Y(_13245_) );
	NAND2X1 NAND2X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_13244_), .B(_13245_), .Y(_13246_) );
	NAND3X1 NAND3X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_13246_), .B(_13233_), .C(_13227_), .Y(_13247_) );
	NAND3X1 NAND3X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_13243_), .B(_13247_), .C(_13242_), .Y(_13248_) );
	AOI21X1 AOI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_13240_), .B(_13248_), .C(_13198_), .Y(_13249_) );
	OAI21X1 OAI21X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_13194_), .B(_13196_), .C(_13172_), .Y(_13251_) );
	NAND3X1 NAND3X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_13193_), .B(_13187_), .C(_13191_), .Y(_13252_) );
	NAND2X1 NAND2X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_13252_), .B(_13251_), .Y(_13253_) );
	NAND3X1 NAND3X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_13243_), .B(_13247_), .C(_13200_), .Y(_13254_) );
	OAI21X1 OAI21X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_13234_), .B(_13238_), .C(_13242_), .Y(_13255_) );
	AOI21X1 AOI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_13255_), .B(_13254_), .C(_13253_), .Y(_13256_) );
	OAI21X1 OAI21X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_13249_), .B(_13256_), .C(_13170_), .Y(_13257_) );
	INVX1 INVX1_1842 ( .gnd(gnd), .vdd(vdd), .A(_12982_), .Y(_13258_) );
	AOI21X1 AOI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_12940_), .B(_12987_), .C(_13258_), .Y(_13259_) );
	NAND3X1 NAND3X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_13254_), .B(_13253_), .C(_13255_), .Y(_13260_) );
	NAND3X1 NAND3X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_13198_), .B(_13248_), .C(_13240_), .Y(_13262_) );
	NAND3X1 NAND3X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_13260_), .B(_13262_), .C(_13259_), .Y(_13263_) );
	AOI21X1 AOI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_13263_), .B(_13257_), .C(_13168_), .Y(_13264_) );
	OAI21X1 OAI21X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_13165_), .B(_13166_), .C(_13122_), .Y(_13265_) );
	NAND3X1 NAND3X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_13157_), .B(_13161_), .C(_13164_), .Y(_13266_) );
	NAND2X1 NAND2X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_13266_), .B(_13265_), .Y(_13267_) );
	NAND3X1 NAND3X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_13260_), .B(_13262_), .C(_13170_), .Y(_13268_) );
	OAI21X1 OAI21X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_13249_), .B(_13256_), .C(_13259_), .Y(_13269_) );
	AOI21X1 AOI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_13269_), .B(_13268_), .C(_13267_), .Y(_13270_) );
	OAI21X1 OAI21X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_13270_), .B(_13264_), .C(_13121_), .Y(_13271_) );
	INVX1 INVX1_1843 ( .gnd(gnd), .vdd(vdd), .A(_12996_), .Y(_13273_) );
	AOI21X1 AOI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_12910_), .B(_13003_), .C(_13273_), .Y(_13274_) );
	NAND3X1 NAND3X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_13268_), .B(_13269_), .C(_13267_), .Y(_13275_) );
	INVX1 INVX1_1844 ( .gnd(gnd), .vdd(vdd), .A(_13268_), .Y(_13276_) );
	AOI21X1 AOI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_13262_), .B(_13260_), .C(_13170_), .Y(_13277_) );
	OAI21X1 OAI21X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(_13276_), .C(_13168_), .Y(_13278_) );
	NAND3X1 NAND3X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_13275_), .B(_13278_), .C(_13274_), .Y(_13279_) );
	AOI21X1 AOI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_13279_), .B(_13271_), .C(_13119_), .Y(_13280_) );
	NAND3X1 NAND3X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_13275_), .B(_13278_), .C(_13121_), .Y(_13281_) );
	OAI21X1 OAI21X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_13270_), .B(_13264_), .C(_13274_), .Y(_13282_) );
	AOI22X1 AOI22X1_296 ( .gnd(gnd), .vdd(vdd), .A(_13113_), .B(_13117_), .C(_13282_), .D(_13281_), .Y(_13284_) );
	OAI21X1 OAI21X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_13284_), .B(_13280_), .C(_13064_), .Y(_13285_) );
	NOR3X1 NOR3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_13016_), .B(_13015_), .C(_13014_), .Y(_13286_) );
	AOI21X1 AOI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_12858_), .B(_13017_), .C(_13286_), .Y(_13287_) );
	NAND3X1 NAND3X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_13108_), .B(_13114_), .C(_13112_), .Y(_13288_) );
	NAND3X1 NAND3X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_13065_), .B(_13116_), .C(_13115_), .Y(_13289_) );
	NAND2X1 NAND2X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_13288_), .B(_13289_), .Y(_13290_) );
	NAND3X1 NAND3X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_13282_), .B(_13290_), .C(_13281_), .Y(_13291_) );
	NAND3X1 NAND3X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_13271_), .B(_13119_), .C(_13279_), .Y(_13292_) );
	NAND3X1 NAND3X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_13291_), .B(_13292_), .C(_13287_), .Y(_13293_) );
	AOI21X1 AOI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_13285_), .B(_13293_), .C(_13062_), .Y(_13295_) );
	NAND3X1 NAND3X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_13291_), .B(_13292_), .C(_13064_), .Y(_13296_) );
	OAI21X1 OAI21X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_13284_), .B(_13280_), .C(_13287_), .Y(_13297_) );
	AOI21X1 AOI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_13297_), .B(_13296_), .C(_13061_), .Y(_13298_) );
	OAI21X1 OAI21X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_13295_), .B(_13298_), .C(_13060_), .Y(_13299_) );
	NAND2X1 NAND2X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_13018_), .B(_13025_), .Y(_13300_) );
	NOR2X1 NOR2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_13028_), .B(_13300_), .Y(_13301_) );
	AOI21X1 AOI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_12800_), .B(_13031_), .C(_13301_), .Y(_13302_) );
	NAND3X1 NAND3X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .B(_13296_), .C(_13297_), .Y(_13303_) );
	NAND3X1 NAND3X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_13062_), .B(_13293_), .C(_13285_), .Y(_13304_) );
	NAND3X1 NAND3X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_13303_), .B(_13304_), .C(_13302_), .Y(_13306_) );
	AOI21X1 AOI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_13306_), .B(_13299_), .C(_13037_), .Y(_13307_) );
	INVX1 INVX1_1845 ( .gnd(gnd), .vdd(vdd), .A(_13037_), .Y(_13308_) );
	NAND3X1 NAND3X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_13303_), .B(_13304_), .C(_13060_), .Y(_13309_) );
	OAI21X1 OAI21X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_13295_), .B(_13298_), .C(_13302_), .Y(_13310_) );
	AOI21X1 AOI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_13309_), .B(_13310_), .C(_13308_), .Y(_13311_) );
	NOR3X1 NOR3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_13307_), .B(_13058_), .C(_13311_), .Y(_13312_) );
	NAND3X1 NAND3X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_13309_), .B(_13310_), .C(_13308_), .Y(_13313_) );
	NAND3X1 NAND3X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_13037_), .B(_13299_), .C(_13306_), .Y(_13314_) );
	AOI21X1 AOI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_13313_), .B(_13314_), .C(_13044_), .Y(_13315_) );
	NOR2X1 NOR2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_13315_), .B(_13312_), .Y(_13317_) );
	XNOR2X1 XNOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_13057_), .B(_13317_), .Y(mulOut_19_) );
	NAND3X1 NAND3X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_13314_), .B(_13313_), .C(_13044_), .Y(_13318_) );
	OAI21X1 OAI21X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_13307_), .B(_13311_), .C(_13058_), .Y(_13319_) );
	AOI22X1 AOI22X1_297 ( .gnd(gnd), .vdd(vdd), .A(_13319_), .B(_13318_), .C(_13048_), .D(_13052_), .Y(_13320_) );
	NAND2X1 NAND2X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_12793_), .B(_13320_), .Y(_13321_) );
	OAI21X1 OAI21X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_13307_), .B(_13311_), .C(_13044_), .Y(_13322_) );
	NAND2X1 NAND2X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_13314_), .B(_13313_), .Y(_13323_) );
	OAI21X1 OAI21X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_13044_), .B(_13323_), .C(_13055_), .Y(_13324_) );
	AOI22X1 AOI22X1_298 ( .gnd(gnd), .vdd(vdd), .A(_13322_), .B(_13324_), .C(_13320_), .D(_12792_), .Y(_13325_) );
	OAI21X1 OAI21X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_13321_), .B(_12331_), .C(_13325_), .Y(_13327_) );
	AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_13304_), .B(_13303_), .Y(_13328_) );
	AOI21X1 AOI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_13291_), .B(_13292_), .C(_13064_), .Y(_13329_) );
	OAI21X1 OAI21X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_13062_), .B(_13329_), .C(_13296_), .Y(_13330_) );
	AOI21X1 AOI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_13278_), .B(_13275_), .C(_13121_), .Y(_13331_) );
	OAI21X1 OAI21X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_13119_), .B(_13331_), .C(_13281_), .Y(_13332_) );
	NAND2X1 NAND2X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_13098_), .B(_13102_), .Y(_13333_) );
	INVX4 INVX4_21 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_20_bF_buf0), .Y(_13334_) );
	NOR2X1 NOR2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf0), .B(_13334_), .Y(_13335_) );
	NAND2X1 NAND2X1_2724 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf1), .B(adder_bOperand_19_bF_buf0), .Y(_13336_) );
	INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_18_bF_buf1), .Y(_13338_) );
	OAI21X1 OAI21X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf0), .B(_13338_), .C(_13066_), .Y(_13339_) );
	OAI21X1 OAI21X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_13068_), .B(_13336_), .C(_13339_), .Y(_13340_) );
	XOR2X1 XOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_13340_), .B(_13335_), .Y(_13341_) );
	OAI21X1 OAI21X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_12806_), .B(_13066_), .C(_13341_), .Y(_13342_) );
	NOR2X1 NOR2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_12806_), .B(_13066_), .Y(_13343_) );
	INVX1 INVX1_1846 ( .gnd(gnd), .vdd(vdd), .A(_13343_), .Y(_13344_) );
	OR2X2 OR2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_13341_), .B(_13344_), .Y(_13345_) );
	AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_13345_), .B(_13342_), .Y(_13346_) );
	INVX1 INVX1_1847 ( .gnd(gnd), .vdd(vdd), .A(_13073_), .Y(_13347_) );
	AOI21X1 AOI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_13083_), .B(_13080_), .C(_13087_), .Y(_13349_) );
	OAI21X1 OAI21X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_13349_), .B(_13347_), .C(_13088_), .Y(_13350_) );
	INVX1 INVX1_1848 ( .gnd(gnd), .vdd(vdd), .A(_13077_), .Y(_13351_) );
	OAI21X1 OAI21X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_12811_), .B(_13351_), .C(_13080_), .Y(_13352_) );
	NAND2X1 NAND2X1_2725 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf0), .B(adder_bOperand_17_bF_buf2), .Y(_13353_) );
	INVX1 INVX1_1849 ( .gnd(gnd), .vdd(vdd), .A(_13353_), .Y(_13354_) );
	AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf2), .B(adder_bOperand_16_bF_buf3), .Y(_13355_) );
	AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf0), .B(adder_bOperand_15_bF_buf1), .Y(_13356_) );
	NAND2X1 NAND2X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_13355_), .B(_13356_), .Y(_13357_) );
	OAI22X1 OAI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf3), .B(_12342_), .C(_12780_), .D(_12131_), .Y(_13358_) );
	NAND3X1 NAND3X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_13354_), .B(_13358_), .C(_13357_), .Y(_13360_) );
	OAI21X1 OAI21X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf2), .B(_12342_), .C(_13356_), .Y(_13361_) );
	OAI21X1 OAI21X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_12131_), .C(_13355_), .Y(_13362_) );
	NAND3X1 NAND3X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_13353_), .B(_13361_), .C(_13362_), .Y(_13363_) );
	NAND2X1 NAND2X1_2727 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf1), .B(adder_bOperand_12_bF_buf0), .Y(_13364_) );
	AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_12864_), .B(_13364_), .Y(_13365_) );
	OAI22X1 OAI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_13084_), .B(_13124_), .C(_13123_), .D(_13365_), .Y(_13366_) );
	NAND3X1 NAND3X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_13360_), .B(_13363_), .C(_13366_), .Y(_13367_) );
	AOI21X1 AOI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_13361_), .B(_13362_), .C(_13353_), .Y(_13368_) );
	AOI21X1 AOI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_13357_), .B(_13358_), .C(_13354_), .Y(_13369_) );
	NOR2X1 NOR2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_12864_), .B(_13364_), .Y(_13371_) );
	AOI21X1 AOI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_13125_), .B(_13150_), .C(_13371_), .Y(_13372_) );
	OAI21X1 OAI21X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_13369_), .B(_13368_), .C(_13372_), .Y(_13373_) );
	NAND3X1 NAND3X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_13352_), .B(_13367_), .C(_13373_), .Y(_13374_) );
	INVX1 INVX1_1850 ( .gnd(gnd), .vdd(vdd), .A(_13352_), .Y(_13375_) );
	NAND3X1 NAND3X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_13360_), .B(_13372_), .C(_13363_), .Y(_13376_) );
	OAI21X1 OAI21X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_13369_), .B(_13368_), .C(_13366_), .Y(_13377_) );
	NAND3X1 NAND3X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_13376_), .B(_13377_), .C(_13375_), .Y(_13378_) );
	NAND3X1 NAND3X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_13374_), .B(_13378_), .C(_13350_), .Y(_13379_) );
	INVX1 INVX1_1851 ( .gnd(gnd), .vdd(vdd), .A(_13088_), .Y(_13380_) );
	AOI21X1 AOI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_13073_), .B(_13093_), .C(_13380_), .Y(_13382_) );
	AOI21X1 AOI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_13377_), .B(_13376_), .C(_13375_), .Y(_13383_) );
	AOI21X1 AOI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_13373_), .B(_13367_), .C(_13352_), .Y(_13384_) );
	OAI21X1 OAI21X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_13383_), .B(_13384_), .C(_13382_), .Y(_13385_) );
	NAND3X1 NAND3X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_13379_), .B(_13385_), .C(_13346_), .Y(_13386_) );
	NAND2X1 NAND2X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_13342_), .B(_13345_), .Y(_13387_) );
	OAI21X1 OAI21X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_13383_), .B(_13384_), .C(_13350_), .Y(_13388_) );
	NAND3X1 NAND3X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_13374_), .B(_13378_), .C(_13382_), .Y(_13389_) );
	NAND3X1 NAND3X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_13387_), .B(_13388_), .C(_13389_), .Y(_13390_) );
	OAI21X1 OAI21X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_13165_), .B(_13164_), .C(_13161_), .Y(_13391_) );
	NAND3X1 NAND3X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_13386_), .B(_13390_), .C(_13391_), .Y(_13393_) );
	AOI21X1 AOI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_13389_), .B(_13388_), .C(_13387_), .Y(_13394_) );
	AOI22X1 AOI22X1_299 ( .gnd(gnd), .vdd(vdd), .A(_13342_), .B(_13345_), .C(_13379_), .D(_13385_), .Y(_13395_) );
	AOI21X1 AOI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_13122_), .B(_13157_), .C(_13166_), .Y(_13396_) );
	OAI21X1 OAI21X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_13395_), .B(_13394_), .C(_13396_), .Y(_13397_) );
	NAND3X1 NAND3X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_13333_), .B(_13397_), .C(_13393_), .Y(_13398_) );
	AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(_13102_), .B(_13098_), .Y(_13399_) );
	NOR3X1 NOR3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_13395_), .B(_13394_), .C(_13396_), .Y(_13400_) );
	AOI21X1 AOI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_13386_), .B(_13390_), .C(_13391_), .Y(_13401_) );
	OAI21X1 OAI21X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(_13400_), .C(_13399_), .Y(_13402_) );
	NAND2X1 NAND2X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_13398_), .B(_13402_), .Y(_13404_) );
	OAI21X1 OAI21X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(_13168_), .C(_13268_), .Y(_13405_) );
	NAND2X1 NAND2X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_13153_), .B(_13158_), .Y(_13406_) );
	NOR2X1 NOR2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf0), .B(_12365_), .Y(_13407_) );
	INVX1 INVX1_1852 ( .gnd(gnd), .vdd(vdd), .A(_13364_), .Y(_13408_) );
	NAND2X1 NAND2X1_2731 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf3), .B(adder_bOperand_13_bF_buf1), .Y(_13409_) );
	INVX1 INVX1_1853 ( .gnd(gnd), .vdd(vdd), .A(_13409_), .Y(_13410_) );
	NAND2X1 NAND2X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_13408_), .B(_13410_), .Y(_13411_) );
	OAI21X1 OAI21X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_17157_), .C(_13124_), .Y(_13412_) );
	NAND3X1 NAND3X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_13407_), .B(_13412_), .C(_13411_), .Y(_13413_) );
	OAI21X1 OAI21X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_13364_), .B(_13409_), .C(_13412_), .Y(_13415_) );
	OAI21X1 OAI21X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf3), .B(_12365_), .C(_13415_), .Y(_13416_) );
	AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_13416_), .B(_13413_), .Y(_13417_) );
	OAI21X1 OAI21X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_13130_), .B(_13146_), .C(_13136_), .Y(_13418_) );
	NAND2X1 NAND2X1_2733 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf4), .B(adder_bOperand_11_bF_buf1), .Y(_13419_) );
	INVX1 INVX1_1854 ( .gnd(gnd), .vdd(vdd), .A(_13419_), .Y(_13420_) );
	AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf2), .B(adder_bOperand_10_bF_buf2), .Y(_13421_) );
	AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf4), .B(aOperand_frameOut_11_bF_buf0), .Y(_13422_) );
	NAND2X1 NAND2X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_13421_), .B(_13422_), .Y(_13423_) );
	NAND2X1 NAND2X1_2735 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf1), .B(adder_bOperand_10_bF_buf1), .Y(_13424_) );
	OAI21X1 OAI21X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf0), .B(_17077_), .C(_13424_), .Y(_13426_) );
	NAND3X1 NAND3X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_13420_), .B(_13426_), .C(_13423_), .Y(_13427_) );
	NAND2X1 NAND2X1_2736 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf3), .B(aOperand_frameOut_11_bF_buf4), .Y(_13428_) );
	NOR2X1 NOR2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_13424_), .B(_13428_), .Y(_13429_) );
	AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_13424_), .B(_13428_), .Y(_13430_) );
	OAI21X1 OAI21X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_13429_), .B(_13430_), .C(_13419_), .Y(_13431_) );
	NAND3X1 NAND3X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_13427_), .B(_13418_), .C(_13431_), .Y(_13432_) );
	AOI21X1 AOI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_13138_), .B(_13135_), .C(_13145_), .Y(_13433_) );
	OAI21X1 OAI21X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_16887_), .C(_13422_), .Y(_13434_) );
	OAI21X1 OAI21X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf3), .B(_17077_), .C(_13421_), .Y(_13435_) );
	AOI21X1 AOI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_13434_), .B(_13435_), .C(_13419_), .Y(_13437_) );
	AOI21X1 AOI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_13423_), .B(_13426_), .C(_13420_), .Y(_13438_) );
	OAI21X1 OAI21X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_13438_), .B(_13437_), .C(_13433_), .Y(_13439_) );
	NAND3X1 NAND3X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_13432_), .B(_13439_), .C(_13417_), .Y(_13440_) );
	NAND2X1 NAND2X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_13413_), .B(_13416_), .Y(_13441_) );
	OAI21X1 OAI21X1_2898 ( .gnd(gnd), .vdd(vdd), .A(_13438_), .B(_13437_), .C(_13418_), .Y(_13442_) );
	NAND3X1 NAND3X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_13427_), .B(_13433_), .C(_13431_), .Y(_13443_) );
	NAND3X1 NAND3X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_13443_), .B(_13442_), .C(_13441_), .Y(_13444_) );
	OAI21X1 OAI21X1_2899 ( .gnd(gnd), .vdd(vdd), .A(_13193_), .B(_13194_), .C(_13191_), .Y(_13445_) );
	AOI21X1 AOI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_13440_), .B(_13444_), .C(_13445_), .Y(_13446_) );
	AOI21X1 AOI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_13442_), .B(_13443_), .C(_13441_), .Y(_13448_) );
	AOI22X1 AOI22X1_300 ( .gnd(gnd), .vdd(vdd), .A(_13413_), .B(_13416_), .C(_13432_), .D(_13439_), .Y(_13449_) );
	AOI21X1 AOI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_13187_), .B(_13172_), .C(_13196_), .Y(_13450_) );
	NOR3X1 NOR3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_13449_), .B(_13448_), .C(_13450_), .Y(_13451_) );
	OAI21X1 OAI21X1_2900 ( .gnd(gnd), .vdd(vdd), .A(_13446_), .B(_13451_), .C(_13406_), .Y(_13452_) );
	INVX1 INVX1_1855 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .Y(_13453_) );
	OAI21X1 OAI21X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_13449_), .B(_13448_), .C(_13450_), .Y(_13454_) );
	NAND3X1 NAND3X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_13444_), .B(_13445_), .C(_13440_), .Y(_13455_) );
	NAND3X1 NAND3X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_13454_), .B(_13455_), .C(_13453_), .Y(_13456_) );
	AOI21X1 AOI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_13243_), .B(_13247_), .C(_13200_), .Y(_13457_) );
	OAI21X1 OAI21X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_13457_), .B(_13198_), .C(_13254_), .Y(_13459_) );
	NAND2X1 NAND2X1_2738 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf1), .B(aOperand_frameOut_13_bF_buf2), .Y(_13460_) );
	OAI21X1 OAI21X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_12924_), .B(_13460_), .C(_13188_), .Y(_13461_) );
	NAND2X1 NAND2X1_2739 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf1), .B(aOperand_frameOut_12_bF_buf3), .Y(_13462_) );
	NAND3X1 NAND3X1_2878 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf1), .B(aOperand_frameOut_14_bF_buf2), .C(_13460_), .Y(_13463_) );
	NAND2X1 NAND2X1_2740 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf0), .B(aOperand_frameOut_14_bF_buf1), .Y(_13464_) );
	NAND3X1 NAND3X1_2879 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf0), .B(aOperand_frameOut_13_bF_buf1), .C(_13464_), .Y(_13465_) );
	AOI21X1 AOI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_13463_), .B(_13465_), .C(_13462_), .Y(_13466_) );
	AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(aOperand_frameOut_14_bF_buf0), .Y(_13467_) );
	NAND2X1 NAND2X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_13180_), .B(_13467_), .Y(_13468_) );
	OAI21X1 OAI21X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf3), .B(_12039_), .C(_13460_), .Y(_13470_) );
	AOI22X1 AOI22X1_301 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf0), .B(aOperand_frameOut_12_bF_buf2), .C(_13470_), .D(_13468_), .Y(_13471_) );
	AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf2), .B(aOperand_frameOut_16_bF_buf2), .Y(_13472_) );
	AOI22X1 AOI22X1_302 ( .gnd(gnd), .vdd(vdd), .A(_12945_), .B(_13472_), .C(_13209_), .D(_13207_), .Y(_13473_) );
	OAI21X1 OAI21X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_13466_), .B(_13471_), .C(_13473_), .Y(_13474_) );
	INVX1 INVX1_1856 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .Y(_13475_) );
	NAND3X1 NAND3X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_13475_), .B(_13470_), .C(_13468_), .Y(_13476_) );
	NAND3X1 NAND3X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_13462_), .B(_13463_), .C(_13465_), .Y(_13477_) );
	NOR2X1 NOR2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_13185_), .B(_13202_), .Y(_13478_) );
	OAI21X1 OAI21X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_13201_), .B(_13478_), .C(_13203_), .Y(_13479_) );
	NAND3X1 NAND3X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .B(_13477_), .C(_13479_), .Y(_13481_) );
	NAND3X1 NAND3X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_13461_), .B(_13474_), .C(_13481_), .Y(_13482_) );
	AOI21X1 AOI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_12918_), .B(_13180_), .C(_13178_), .Y(_13483_) );
	AOI21X1 AOI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_13476_), .B(_13477_), .C(_13479_), .Y(_13484_) );
	NOR3X1 NOR3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_13473_), .B(_13466_), .C(_13471_), .Y(_13485_) );
	OAI21X1 OAI21X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .B(_13485_), .C(_13483_), .Y(_13486_) );
	NAND2X1 NAND2X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_13482_), .B(_13486_), .Y(_13487_) );
	AOI21X1 AOI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .B(_13232_), .C(_13214_), .Y(_13488_) );
	OAI21X1 OAI21X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_13246_), .B(_13488_), .C(_13236_), .Y(_13489_) );
	NAND2X1 NAND2X1_2743 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf0), .B(aOperand_frameOut_15_bF_buf2), .Y(_13490_) );
	AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf2), .B(aOperand_frameOut_17_bF_buf3), .Y(_13492_) );
	NAND2X1 NAND2X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_13472_), .B(_13492_), .Y(_13493_) );
	NAND2X1 NAND2X1_2745 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf1), .B(aOperand_frameOut_16_bF_buf1), .Y(_13494_) );
	NAND2X1 NAND2X1_2746 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf1), .B(aOperand_frameOut_17_bF_buf2), .Y(_13495_) );
	NAND2X1 NAND2X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13495_), .Y(_13496_) );
	NAND3X1 NAND3X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .B(_13496_), .C(_13493_), .Y(_13497_) );
	INVX1 INVX1_1857 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .Y(_13498_) );
	OAI21X1 OAI21X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_12461_), .C(_13492_), .Y(_13499_) );
	OAI21X1 OAI21X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf3), .B(_12708_), .C(_13472_), .Y(_13500_) );
	NAND3X1 NAND3X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .B(_13499_), .C(_13500_), .Y(_13501_) );
	AOI22X1 AOI22X1_303 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .B(aOperand_frameOut_19_bF_buf1), .C(adder_bOperand_1_bF_buf1), .D(aOperand_frameOut_18_bF_buf4), .Y(_13503_) );
	OAI21X1 OAI21X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_13215_), .B(_13503_), .C(_13223_), .Y(_13504_) );
	NAND2X1 NAND2X1_2748 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf3), .B(aOperand_frameOut_18_bF_buf3), .Y(_13505_) );
	NAND2X1 NAND2X1_2749 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf0), .B(aOperand_frameOut_19_bF_buf0), .Y(_13506_) );
	NAND3X1 NAND3X1_2886 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_20_bF_buf1), .C(_13506_), .Y(_13507_) );
	NAND2X1 NAND2X1_2750 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_20_bF_buf0), .Y(_13508_) );
	NAND3X1 NAND3X1_2887 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf6), .B(aOperand_frameOut_19_bF_buf4), .C(_13508_), .Y(_13509_) );
	AOI21X1 AOI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_13507_), .B(_13509_), .C(_13505_), .Y(_13510_) );
	AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(aOperand_frameOut_20_bF_buf4), .Y(_13511_) );
	NAND2X1 NAND2X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_13222_), .B(_13511_), .Y(_13512_) );
	INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_20_bF_buf3), .Y(_13514_) );
	OAI21X1 OAI21X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf2), .B(_13514_), .C(_13506_), .Y(_13515_) );
	AOI22X1 AOI22X1_304 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf2), .B(aOperand_frameOut_18_bF_buf2), .C(_13515_), .D(_13512_), .Y(_13516_) );
	OAI21X1 OAI21X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_13510_), .B(_13516_), .C(_13504_), .Y(_13517_) );
	INVX1 INVX1_1858 ( .gnd(gnd), .vdd(vdd), .A(_12962_), .Y(_13518_) );
	INVX1 INVX1_1859 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .Y(_13519_) );
	AOI22X1 AOI22X1_305 ( .gnd(gnd), .vdd(vdd), .A(_13518_), .B(_13519_), .C(_13230_), .D(_13225_), .Y(_13520_) );
	INVX1 INVX1_1860 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .Y(_13521_) );
	NAND3X1 NAND3X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_13521_), .B(_13515_), .C(_13512_), .Y(_13522_) );
	NAND3X1 NAND3X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .B(_13507_), .C(_13509_), .Y(_13523_) );
	NAND3X1 NAND3X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_13523_), .B(_13520_), .C(_13522_), .Y(_13525_) );
	AOI22X1 AOI22X1_306 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13501_), .C(_13525_), .D(_13517_), .Y(_13526_) );
	NAND3X1 NAND3X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_13498_), .B(_13496_), .C(_13493_), .Y(_13527_) );
	NAND3X1 NAND3X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_13490_), .B(_13499_), .C(_13500_), .Y(_13528_) );
	NAND3X1 NAND3X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_13523_), .B(_13504_), .C(_13522_), .Y(_13529_) );
	OAI21X1 OAI21X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_13510_), .B(_13516_), .C(_13520_), .Y(_13530_) );
	AOI22X1 AOI22X1_307 ( .gnd(gnd), .vdd(vdd), .A(_13527_), .B(_13528_), .C(_13529_), .D(_13530_), .Y(_13531_) );
	OAI21X1 OAI21X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13531_), .C(_13489_), .Y(_13532_) );
	NOR3X1 NOR3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_13229_), .B(_13221_), .C(_13226_), .Y(_13533_) );
	AOI21X1 AOI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_13235_), .B(_13237_), .C(_13533_), .Y(_13534_) );
	NAND2X1 NAND2X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13501_), .Y(_13536_) );
	NAND3X1 NAND3X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .B(_13529_), .C(_13530_), .Y(_13537_) );
	NAND2X1 NAND2X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_13527_), .B(_13528_), .Y(_13538_) );
	NAND3X1 NAND3X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_13525_), .B(_13538_), .C(_13517_), .Y(_13539_) );
	NAND3X1 NAND3X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_13537_), .B(_13539_), .C(_13534_), .Y(_13540_) );
	AOI21X1 AOI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_13532_), .B(_13540_), .C(_13487_), .Y(_13541_) );
	OAI21X1 OAI21X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_13484_), .B(_13485_), .C(_13461_), .Y(_13542_) );
	NAND3X1 NAND3X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_13483_), .B(_13474_), .C(_13481_), .Y(_13543_) );
	NAND2X1 NAND2X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_13543_), .B(_13542_), .Y(_13544_) );
	NAND3X1 NAND3X1_2898 ( .gnd(gnd), .vdd(vdd), .A(_13537_), .B(_13539_), .C(_13489_), .Y(_13545_) );
	OAI21X1 OAI21X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13531_), .C(_13534_), .Y(_13547_) );
	AOI21X1 AOI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_13547_), .B(_13545_), .C(_13544_), .Y(_13548_) );
	OAI21X1 OAI21X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_13541_), .B(_13548_), .C(_13459_), .Y(_13549_) );
	INVX1 INVX1_1861 ( .gnd(gnd), .vdd(vdd), .A(_13254_), .Y(_13550_) );
	AOI21X1 AOI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_13253_), .B(_13255_), .C(_13550_), .Y(_13551_) );
	NAND3X1 NAND3X1_2899 ( .gnd(gnd), .vdd(vdd), .A(_13545_), .B(_13544_), .C(_13547_), .Y(_13552_) );
	NAND3X1 NAND3X1_2900 ( .gnd(gnd), .vdd(vdd), .A(_13487_), .B(_13540_), .C(_13532_), .Y(_13553_) );
	NAND3X1 NAND3X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_13552_), .B(_13553_), .C(_13551_), .Y(_13554_) );
	AOI22X1 AOI22X1_308 ( .gnd(gnd), .vdd(vdd), .A(_13452_), .B(_13456_), .C(_13549_), .D(_13554_), .Y(_13555_) );
	NAND3X1 NAND3X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .B(_13455_), .C(_13454_), .Y(_13556_) );
	OAI21X1 OAI21X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_13446_), .B(_13451_), .C(_13453_), .Y(_13558_) );
	NAND3X1 NAND3X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_13552_), .B(_13553_), .C(_13459_), .Y(_13559_) );
	OAI21X1 OAI21X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_13541_), .B(_13548_), .C(_13551_), .Y(_13560_) );
	AOI22X1 AOI22X1_309 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_13558_), .C(_13559_), .D(_13560_), .Y(_13561_) );
	OAI21X1 OAI21X1_2921 ( .gnd(gnd), .vdd(vdd), .A(_13561_), .B(_13555_), .C(_13405_), .Y(_13562_) );
	AOI21X1 AOI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_13267_), .B(_13269_), .C(_13276_), .Y(_13563_) );
	NAND2X1 NAND2X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_13456_), .B(_13452_), .Y(_13564_) );
	NAND3X1 NAND3X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_13559_), .B(_13560_), .C(_13564_), .Y(_13565_) );
	NAND2X1 NAND2X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_13558_), .Y(_13566_) );
	INVX1 INVX1_1862 ( .gnd(gnd), .vdd(vdd), .A(_13559_), .Y(_13567_) );
	AOI21X1 AOI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_13553_), .B(_13552_), .C(_13459_), .Y(_13569_) );
	OAI21X1 OAI21X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_13569_), .B(_13567_), .C(_13566_), .Y(_13570_) );
	NAND3X1 NAND3X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_13565_), .B(_13563_), .C(_13570_), .Y(_13571_) );
	AOI21X1 AOI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_13571_), .B(_13562_), .C(_13404_), .Y(_13572_) );
	OAI21X1 OAI21X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(_13400_), .C(_13333_), .Y(_13573_) );
	NAND3X1 NAND3X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .B(_13393_), .C(_13399_), .Y(_13574_) );
	NAND2X1 NAND2X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_13574_), .B(_13573_), .Y(_13575_) );
	NAND3X1 NAND3X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_13405_), .B(_13565_), .C(_13570_), .Y(_13576_) );
	OAI21X1 OAI21X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_13561_), .B(_13555_), .C(_13563_), .Y(_13577_) );
	AOI21X1 AOI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_13576_), .B(_13577_), .C(_13575_), .Y(_13578_) );
	OAI21X1 OAI21X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .B(_13578_), .C(_13332_), .Y(_13580_) );
	NOR3X1 NOR3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_13270_), .B(_13264_), .C(_13274_), .Y(_13581_) );
	AOI21X1 AOI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_13290_), .B(_13282_), .C(_13581_), .Y(_13582_) );
	NAND3X1 NAND3X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_13577_), .B(_13576_), .C(_13575_), .Y(_13583_) );
	NOR3X1 NOR3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_13561_), .B(_13555_), .C(_13563_), .Y(_13584_) );
	AOI21X1 AOI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13565_), .C(_13405_), .Y(_13585_) );
	OAI21X1 OAI21X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_13585_), .B(_13584_), .C(_13404_), .Y(_13586_) );
	NAND3X1 NAND3X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .B(_13586_), .C(_13582_), .Y(_13587_) );
	AOI22X1 AOI22X1_310 ( .gnd(gnd), .vdd(vdd), .A(_13108_), .B(_13113_), .C(_13580_), .D(_13587_), .Y(_13588_) );
	NAND2X1 NAND2X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_13108_), .B(_13113_), .Y(_13589_) );
	NAND3X1 NAND3X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .B(_13332_), .C(_13586_), .Y(_13590_) );
	OAI21X1 OAI21X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_13572_), .B(_13578_), .C(_13582_), .Y(_13591_) );
	AOI21X1 AOI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_13590_), .B(_13591_), .C(_13589_), .Y(_13592_) );
	OAI21X1 OAI21X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_13588_), .B(_13592_), .C(_13330_), .Y(_13593_) );
	NOR3X1 NOR3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_13284_), .B(_13280_), .C(_13287_), .Y(_13594_) );
	AOI21X1 AOI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .B(_13297_), .C(_13594_), .Y(_13595_) );
	NAND3X1 NAND3X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .B(_13591_), .C(_13590_), .Y(_13596_) );
	INVX1 INVX1_1863 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .Y(_13597_) );
	NAND3X1 NAND3X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_13597_), .B(_13580_), .C(_13587_), .Y(_13598_) );
	NAND3X1 NAND3X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_13596_), .B(_13598_), .C(_13595_), .Y(_13599_) );
	AOI22X1 AOI22X1_311 ( .gnd(gnd), .vdd(vdd), .A(_13060_), .B(_13328_), .C(_13593_), .D(_13599_), .Y(_13602_) );
	NAND3X1 NAND3X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_13596_), .B(_13598_), .C(_13330_), .Y(_13603_) );
	OAI21X1 OAI21X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_13588_), .B(_13592_), .C(_13595_), .Y(_13604_) );
	AOI21X1 AOI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_13604_), .B(_13603_), .C(_13309_), .Y(_13605_) );
	OAI21X1 OAI21X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_13602_), .B(_13605_), .C(_13307_), .Y(_13606_) );
	AOI21X1 AOI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_13599_), .B(_13593_), .C(_13309_), .Y(_13607_) );
	AOI22X1 AOI22X1_312 ( .gnd(gnd), .vdd(vdd), .A(_13328_), .B(_13060_), .C(_13603_), .D(_13604_), .Y(_13608_) );
	OAI21X1 OAI21X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_13608_), .B(_13607_), .C(_13313_), .Y(_13609_) );
	NAND2X1 NAND2X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_13606_), .B(_13609_), .Y(_13610_) );
	XNOR2X1 XNOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_13327_), .B(_13610_), .Y(mulOut_20_) );
	NOR3X1 NOR3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_13608_), .B(_13607_), .C(_13313_), .Y(_13611_) );
	AOI21X1 AOI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_13327_), .B(_13609_), .C(_13611_), .Y(_13612_) );
	INVX1 INVX1_1864 ( .gnd(gnd), .vdd(vdd), .A(_13607_), .Y(_13613_) );
	INVX1 INVX1_1865 ( .gnd(gnd), .vdd(vdd), .A(_13603_), .Y(_13614_) );
	NAND2X1 NAND2X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_13590_), .B(_13596_), .Y(_13615_) );
	INVX1 INVX1_1866 ( .gnd(gnd), .vdd(vdd), .A(_13345_), .Y(_13616_) );
	OAI21X1 OAI21X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_13401_), .B(_13399_), .C(_13393_), .Y(_13617_) );
	NAND2X1 NAND2X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_13616_), .B(_13617_), .Y(_13618_) );
	INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .Y(_13619_) );
	NOR2X1 NOR2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_13616_), .B(_13617_), .Y(_13620_) );
	NOR2X1 NOR2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_13620_), .B(_13619_), .Y(_13623_) );
	OAI21X1 OAI21X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_13404_), .B(_13585_), .C(_13576_), .Y(_13624_) );
	AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_13386_), .B(_13379_), .Y(_13625_) );
	NAND2X1 NAND2X1_2762 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf4), .B(adder_bOperand_21_bF_buf3), .Y(_13626_) );
	NAND2X1 NAND2X1_2763 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf0), .B(adder_bOperand_18_bF_buf0), .Y(_13627_) );
	NOR2X1 NOR2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_13066_), .B(_13627_), .Y(_13628_) );
	AOI21X1 AOI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_13339_), .B(_13335_), .C(_13628_), .Y(_13629_) );
	INVX1 INVX1_1867 ( .gnd(gnd), .vdd(vdd), .A(_13629_), .Y(_13630_) );
	NOR2X1 NOR2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_13334_), .Y(_13631_) );
	INVX1 INVX1_1868 ( .gnd(gnd), .vdd(vdd), .A(_13631_), .Y(_13632_) );
	NAND2X1 NAND2X1_2764 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf4), .B(adder_bOperand_19_bF_buf3), .Y(_13634_) );
	OAI21X1 OAI21X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_13338_), .C(_13336_), .Y(_13635_) );
	OAI21X1 OAI21X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_13627_), .B(_13634_), .C(_13635_), .Y(_13636_) );
	OR2X2 OR2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_13636_), .B(_13632_), .Y(_13637_) );
	OAI21X1 OAI21X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_13334_), .C(_13636_), .Y(_13638_) );
	AOI21X1 AOI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_13637_), .B(_13638_), .C(_13630_), .Y(_13639_) );
	NOR2X1 NOR2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_13632_), .B(_13636_), .Y(_13640_) );
	INVX1 INVX1_1869 ( .gnd(gnd), .vdd(vdd), .A(_13627_), .Y(_13641_) );
	INVX1 INVX1_1870 ( .gnd(gnd), .vdd(vdd), .A(_13634_), .Y(_13642_) );
	NAND2X1 NAND2X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_13641_), .B(_13642_), .Y(_13643_) );
	AOI21X1 AOI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_13643_), .B(_13635_), .C(_13631_), .Y(_13645_) );
	NOR3X1 NOR3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_13629_), .B(_13645_), .C(_13640_), .Y(_13646_) );
	OAI21X1 OAI21X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_13646_), .B(_13639_), .C(_13626_), .Y(_13647_) );
	INVX1 INVX1_1871 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .Y(_13648_) );
	OAI21X1 OAI21X1_2938 ( .gnd(gnd), .vdd(vdd), .A(_13645_), .B(_13640_), .C(_13629_), .Y(_13649_) );
	NAND3X1 NAND3X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_13638_), .B(_13630_), .C(_13637_), .Y(_13650_) );
	NAND3X1 NAND3X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_13648_), .B(_13649_), .C(_13650_), .Y(_13651_) );
	AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13651_), .Y(_13652_) );
	NAND2X1 NAND2X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_13367_), .B(_13374_), .Y(_13653_) );
	NAND2X1 NAND2X1_2767 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf4), .B(adder_bOperand_16_bF_buf2), .Y(_13654_) );
	OAI21X1 OAI21X1_2939 ( .gnd(gnd), .vdd(vdd), .A(_13351_), .B(_13654_), .C(_13360_), .Y(_13656_) );
	NAND2X1 NAND2X1_2768 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf1), .B(adder_bOperand_17_bF_buf1), .Y(_13657_) );
	INVX1 INVX1_1872 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .Y(_13658_) );
	AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf2), .B(adder_bOperand_16_bF_buf1), .Y(_13659_) );
	NAND2X1 NAND2X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .B(_13659_), .Y(_13660_) );
	OAI21X1 OAI21X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf2), .B(_12131_), .C(_13654_), .Y(_13661_) );
	NAND3X1 NAND3X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_13658_), .B(_13661_), .C(_13660_), .Y(_13662_) );
	NAND2X1 NAND2X1_2770 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf1), .B(adder_bOperand_15_bF_buf0), .Y(_13663_) );
	NOR2X1 NOR2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_13654_), .B(_13663_), .Y(_13664_) );
	AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_13654_), .B(_13663_), .Y(_13665_) );
	OAI21X1 OAI21X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_13664_), .B(_13665_), .C(_13657_), .Y(_13667_) );
	AOI22X1 AOI22X1_313 ( .gnd(gnd), .vdd(vdd), .A(_13408_), .B(_13410_), .C(_13407_), .D(_13412_), .Y(_13668_) );
	INVX1 INVX1_1873 ( .gnd(gnd), .vdd(vdd), .A(_13668_), .Y(_13669_) );
	NAND3X1 NAND3X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_13662_), .B(_13667_), .C(_13669_), .Y(_13670_) );
	INVX1 INVX1_1874 ( .gnd(gnd), .vdd(vdd), .A(_13662_), .Y(_13671_) );
	AOI21X1 AOI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_13660_), .B(_13661_), .C(_13658_), .Y(_13672_) );
	OAI21X1 OAI21X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_13672_), .B(_13671_), .C(_13668_), .Y(_13673_) );
	NAND3X1 NAND3X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_13656_), .B(_13670_), .C(_13673_), .Y(_13674_) );
	INVX1 INVX1_1875 ( .gnd(gnd), .vdd(vdd), .A(_13656_), .Y(_13675_) );
	NAND2X1 NAND2X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_13662_), .B(_13667_), .Y(_13676_) );
	NOR2X1 NOR2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_13668_), .B(_13676_), .Y(_13678_) );
	AOI21X1 AOI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_13667_), .B(_13662_), .C(_13669_), .Y(_13679_) );
	OAI21X1 OAI21X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_13679_), .B(_13678_), .C(_13675_), .Y(_13680_) );
	NAND3X1 NAND3X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(_13680_), .C(_13653_), .Y(_13681_) );
	INVX1 INVX1_1876 ( .gnd(gnd), .vdd(vdd), .A(_13367_), .Y(_13682_) );
	AOI21X1 AOI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_13352_), .B(_13373_), .C(_13682_), .Y(_13683_) );
	NAND3X1 NAND3X1_2921 ( .gnd(gnd), .vdd(vdd), .A(_13662_), .B(_13668_), .C(_13667_), .Y(_13684_) );
	OAI21X1 OAI21X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_13672_), .B(_13671_), .C(_13669_), .Y(_13685_) );
	AOI21X1 AOI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_13685_), .B(_13684_), .C(_13675_), .Y(_13686_) );
	AOI21X1 AOI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_13673_), .B(_13670_), .C(_13656_), .Y(_13687_) );
	OAI21X1 OAI21X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_13686_), .B(_13687_), .C(_13683_), .Y(_13689_) );
	NAND3X1 NAND3X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_13681_), .B(_13689_), .C(_13652_), .Y(_13690_) );
	NAND2X1 NAND2X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_13651_), .B(_13647_), .Y(_13691_) );
	OAI21X1 OAI21X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_13686_), .B(_13687_), .C(_13653_), .Y(_13692_) );
	NAND3X1 NAND3X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_13674_), .B(_13683_), .C(_13680_), .Y(_13693_) );
	NAND3X1 NAND3X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_13693_), .B(_13691_), .C(_13692_), .Y(_13694_) );
	OAI21X1 OAI21X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_13446_), .B(_13453_), .C(_13455_), .Y(_13695_) );
	NAND3X1 NAND3X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .B(_13695_), .C(_13690_), .Y(_13696_) );
	AOI21X1 AOI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_13692_), .B(_13693_), .C(_13691_), .Y(_13697_) );
	AOI22X1 AOI22X1_314 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13651_), .C(_13681_), .D(_13689_), .Y(_13698_) );
	AOI21X1 AOI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .B(_13454_), .C(_13451_), .Y(_13700_) );
	OAI21X1 OAI21X1_2948 ( .gnd(gnd), .vdd(vdd), .A(_13698_), .B(_13697_), .C(_13700_), .Y(_13701_) );
	NAND3X1 NAND3X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_13625_), .B(_13696_), .C(_13701_), .Y(_13702_) );
	NAND2X1 NAND2X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_13379_), .B(_13386_), .Y(_13703_) );
	NAND3X1 NAND3X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_13694_), .B(_13700_), .C(_13690_), .Y(_13704_) );
	OAI21X1 OAI21X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_13698_), .B(_13697_), .C(_13695_), .Y(_13705_) );
	NAND3X1 NAND3X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_13703_), .B(_13704_), .C(_13705_), .Y(_13706_) );
	NAND2X1 NAND2X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_13702_), .B(_13706_), .Y(_13707_) );
	OAI21X1 OAI21X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_13569_), .B(_13566_), .C(_13559_), .Y(_13708_) );
	NAND2X1 NAND2X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_13432_), .B(_13440_), .Y(_13709_) );
	NOR2X1 NOR2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_12365_), .Y(_13711_) );
	NAND2X1 NAND2X1_2776 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf3), .B(adder_bOperand_12_bF_buf3), .Y(_13712_) );
	NOR2X1 NOR2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_13409_), .B(_13712_), .Y(_13713_) );
	INVX1 INVX1_1877 ( .gnd(gnd), .vdd(vdd), .A(_13713_), .Y(_13714_) );
	OAI21X1 OAI21X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf0), .B(_17157_), .C(_13409_), .Y(_13715_) );
	NAND3X1 NAND3X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_13711_), .B(_13715_), .C(_13714_), .Y(_13716_) );
	INVX1 INVX1_1878 ( .gnd(gnd), .vdd(vdd), .A(_13711_), .Y(_13717_) );
	INVX1 INVX1_1879 ( .gnd(gnd), .vdd(vdd), .A(_13715_), .Y(_13718_) );
	OAI21X1 OAI21X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_13713_), .B(_13718_), .C(_13717_), .Y(_13719_) );
	AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_13719_), .B(_13716_), .Y(_13720_) );
	OAI21X1 OAI21X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_13419_), .B(_13430_), .C(_13423_), .Y(_13722_) );
	NAND2X1 NAND2X1_2777 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf0), .B(adder_bOperand_11_bF_buf0), .Y(_13723_) );
	INVX1 INVX1_1880 ( .gnd(gnd), .vdd(vdd), .A(_13723_), .Y(_13724_) );
	AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf0), .B(aOperand_frameOut_11_bF_buf3), .Y(_13725_) );
	AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf2), .B(aOperand_frameOut_12_bF_buf1), .Y(_13726_) );
	NAND2X1 NAND2X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_13725_), .B(_13726_), .Y(_13727_) );
	NAND2X1 NAND2X1_2779 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf4), .B(aOperand_frameOut_11_bF_buf2), .Y(_13728_) );
	OAI21X1 OAI21X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf2), .B(_17236__bF_buf1), .C(_13728_), .Y(_13729_) );
	NAND3X1 NAND3X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_13724_), .B(_13729_), .C(_13727_), .Y(_13730_) );
	NAND2X1 NAND2X1_2780 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf1), .B(aOperand_frameOut_12_bF_buf0), .Y(_13731_) );
	NOR2X1 NOR2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_13728_), .B(_13731_), .Y(_13732_) );
	NOR2X1 NOR2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_13725_), .B(_13726_), .Y(_13733_) );
	OAI21X1 OAI21X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_13732_), .B(_13733_), .C(_13723_), .Y(_13734_) );
	NAND3X1 NAND3X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_13722_), .B(_13730_), .C(_13734_), .Y(_13735_) );
	AOI21X1 AOI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_13426_), .B(_13420_), .C(_13429_), .Y(_13736_) );
	OAI21X1 OAI21X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_16887_), .B(_17077_), .C(_13726_), .Y(_13737_) );
	OAI21X1 OAI21X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf1), .B(_17236__bF_buf0), .C(_13725_), .Y(_13738_) );
	AOI21X1 AOI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_13737_), .B(_13738_), .C(_13723_), .Y(_13739_) );
	AOI21X1 AOI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_13727_), .B(_13729_), .C(_13724_), .Y(_13740_) );
	OAI21X1 OAI21X1_2958 ( .gnd(gnd), .vdd(vdd), .A(_13740_), .B(_13739_), .C(_13736_), .Y(_13741_) );
	NAND3X1 NAND3X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_13735_), .B(_13741_), .C(_13720_), .Y(_13743_) );
	NAND2X1 NAND2X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_13716_), .B(_13719_), .Y(_13744_) );
	OAI21X1 OAI21X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_13740_), .B(_13739_), .C(_13722_), .Y(_13745_) );
	NAND3X1 NAND3X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_13730_), .B(_13736_), .C(_13734_), .Y(_13746_) );
	NAND3X1 NAND3X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_13746_), .B(_13745_), .C(_13744_), .Y(_13747_) );
	OAI21X1 OAI21X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_13483_), .B(_13484_), .C(_13481_), .Y(_13748_) );
	AOI21X1 AOI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_13743_), .B(_13747_), .C(_13748_), .Y(_13749_) );
	AOI21X1 AOI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_13745_), .B(_13746_), .C(_13744_), .Y(_13750_) );
	AOI22X1 AOI22X1_315 ( .gnd(gnd), .vdd(vdd), .A(_13716_), .B(_13719_), .C(_13735_), .D(_13741_), .Y(_13751_) );
	AOI21X1 AOI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_13461_), .B(_13474_), .C(_13485_), .Y(_13752_) );
	NOR3X1 NOR3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_13751_), .B(_13750_), .C(_13752_), .Y(_13754_) );
	OAI21X1 OAI21X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_13749_), .B(_13754_), .C(_13709_), .Y(_13755_) );
	INVX1 INVX1_1881 ( .gnd(gnd), .vdd(vdd), .A(_13709_), .Y(_13756_) );
	OAI21X1 OAI21X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_13751_), .B(_13750_), .C(_13752_), .Y(_13757_) );
	NAND3X1 NAND3X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_13747_), .B(_13748_), .C(_13743_), .Y(_13758_) );
	NAND3X1 NAND3X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_13758_), .B(_13757_), .C(_13756_), .Y(_13759_) );
	NAND2X1 NAND2X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_13759_), .B(_13755_), .Y(_13760_) );
	AOI21X1 AOI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_13537_), .B(_13539_), .C(_13489_), .Y(_13761_) );
	OAI21X1 OAI21X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_13761_), .B(_13487_), .C(_13545_), .Y(_13762_) );
	NAND2X1 NAND2X1_2783 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(aOperand_frameOut_14_bF_buf4), .Y(_13763_) );
	OAI21X1 OAI21X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_13176_), .B(_13763_), .C(_13476_), .Y(_13765_) );
	NAND2X1 NAND2X1_2784 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf4), .B(aOperand_frameOut_13_bF_buf0), .Y(_13766_) );
	INVX1 INVX1_1882 ( .gnd(gnd), .vdd(vdd), .A(_13766_), .Y(_13767_) );
	AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf4), .B(aOperand_frameOut_15_bF_buf1), .Y(_13768_) );
	NAND2X1 NAND2X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_13467_), .B(_13768_), .Y(_13769_) );
	OAI21X1 OAI21X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf2), .B(_12233_), .C(_13763_), .Y(_13770_) );
	NAND3X1 NAND3X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_13767_), .B(_13770_), .C(_13769_), .Y(_13771_) );
	NAND3X1 NAND3X1_2938 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf4), .B(aOperand_frameOut_15_bF_buf0), .C(_13763_), .Y(_13772_) );
	NAND2X1 NAND2X1_2786 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf3), .B(aOperand_frameOut_15_bF_buf4), .Y(_13773_) );
	NAND3X1 NAND3X1_2939 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf3), .B(aOperand_frameOut_14_bF_buf3), .C(_13773_), .Y(_13774_) );
	NAND3X1 NAND3X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_13766_), .B(_13772_), .C(_13774_), .Y(_13776_) );
	AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf0), .B(aOperand_frameOut_17_bF_buf1), .Y(_13777_) );
	AOI22X1 AOI22X1_316 ( .gnd(gnd), .vdd(vdd), .A(_13202_), .B(_13777_), .C(_13498_), .D(_13496_), .Y(_13778_) );
	INVX1 INVX1_1883 ( .gnd(gnd), .vdd(vdd), .A(_13778_), .Y(_13779_) );
	AOI21X1 AOI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_13771_), .B(_13776_), .C(_13779_), .Y(_13780_) );
	AOI21X1 AOI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_13772_), .B(_13774_), .C(_13766_), .Y(_13781_) );
	AOI21X1 AOI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_13769_), .B(_13770_), .C(_13767_), .Y(_13782_) );
	NOR3X1 NOR3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_13778_), .B(_13781_), .C(_13782_), .Y(_13783_) );
	OAI21X1 OAI21X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_13780_), .B(_13783_), .C(_13765_), .Y(_13784_) );
	INVX1 INVX1_1884 ( .gnd(gnd), .vdd(vdd), .A(_13765_), .Y(_13785_) );
	OAI21X1 OAI21X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_13781_), .B(_13782_), .C(_13778_), .Y(_13787_) );
	NAND3X1 NAND3X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_13771_), .B(_13776_), .C(_13779_), .Y(_13788_) );
	NAND3X1 NAND3X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_13787_), .B(_13788_), .C(_13785_), .Y(_13789_) );
	NAND2X1 NAND2X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_13789_), .B(_13784_), .Y(_13790_) );
	AOI21X1 AOI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_13522_), .B(_13523_), .C(_13504_), .Y(_13791_) );
	OAI21X1 OAI21X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_13538_), .B(_13791_), .C(_13529_), .Y(_13792_) );
	NAND2X1 NAND2X1_2788 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf4), .B(aOperand_frameOut_16_bF_buf0), .Y(_13793_) );
	AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf0), .B(aOperand_frameOut_18_bF_buf1), .Y(_13794_) );
	NAND2X1 NAND2X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_13777_), .B(_13794_), .Y(_13795_) );
	INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_18_bF_buf0), .Y(_13796_) );
	OAI22X1 OAI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf2), .B(_13796_), .C(_12266_), .D(_12708_), .Y(_13798_) );
	NAND3X1 NAND3X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_13793_), .B(_13798_), .C(_13795_), .Y(_13799_) );
	INVX1 INVX1_1885 ( .gnd(gnd), .vdd(vdd), .A(_13793_), .Y(_13800_) );
	OAI21X1 OAI21X1_2969 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_12708_), .C(_13794_), .Y(_13801_) );
	OAI21X1 OAI21X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf1), .B(_13796_), .C(_13777_), .Y(_13802_) );
	NAND3X1 NAND3X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_13800_), .B(_13801_), .C(_13802_), .Y(_13803_) );
	NAND2X1 NAND2X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_13799_), .B(_13803_), .Y(_13804_) );
	AOI22X1 AOI22X1_317 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_20_bF_buf2), .C(adder_bOperand_1_bF_buf4), .D(aOperand_frameOut_19_bF_buf3), .Y(_13805_) );
	OAI21X1 OAI21X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .B(_13805_), .C(_13512_), .Y(_13806_) );
	NAND2X1 NAND2X1_2791 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf1), .B(aOperand_frameOut_19_bF_buf2), .Y(_13807_) );
	INVX1 INVX1_1886 ( .gnd(gnd), .vdd(vdd), .A(_13807_), .Y(_13809_) );
	AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(aOperand_frameOut_21_bF_buf4), .Y(_13810_) );
	NAND2X1 NAND2X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_13511_), .B(_13810_), .Y(_13811_) );
	INVX4 INVX4_22 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_21_bF_buf3), .Y(_13812_) );
	NAND2X1 NAND2X1_2793 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf3), .B(aOperand_frameOut_20_bF_buf1), .Y(_13813_) );
	OAI21X1 OAI21X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf1), .B(_13812_), .C(_13813_), .Y(_13814_) );
	NAND3X1 NAND3X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_13809_), .B(_13814_), .C(_13811_), .Y(_13815_) );
	NAND2X1 NAND2X1_2794 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .B(aOperand_frameOut_21_bF_buf2), .Y(_13816_) );
	NOR2X1 NOR2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_13813_), .B(_13816_), .Y(_13817_) );
	AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_13813_), .B(_13816_), .Y(_13818_) );
	OAI21X1 OAI21X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_13817_), .B(_13818_), .C(_13807_), .Y(_13820_) );
	NAND3X1 NAND3X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_13806_), .B(_13815_), .C(_13820_), .Y(_13821_) );
	AOI22X1 AOI22X1_318 ( .gnd(gnd), .vdd(vdd), .A(_13222_), .B(_13511_), .C(_13521_), .D(_13515_), .Y(_13822_) );
	NAND3X1 NAND3X1_2947 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(aOperand_frameOut_21_bF_buf1), .C(_13813_), .Y(_13823_) );
	NAND3X1 NAND3X1_2948 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .B(aOperand_frameOut_20_bF_buf0), .C(_13816_), .Y(_13824_) );
	AOI21X1 AOI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_13823_), .B(_13824_), .C(_13807_), .Y(_13825_) );
	AOI22X1 AOI22X1_319 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf0), .B(aOperand_frameOut_19_bF_buf1), .C(_13814_), .D(_13811_), .Y(_13826_) );
	OAI21X1 OAI21X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_13825_), .B(_13826_), .C(_13822_), .Y(_13827_) );
	NAND3X1 NAND3X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_13804_), .B(_13821_), .C(_13827_), .Y(_13828_) );
	AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_13803_), .B(_13799_), .Y(_13829_) );
	OAI21X1 OAI21X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_13825_), .B(_13826_), .C(_13806_), .Y(_13831_) );
	NAND3X1 NAND3X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_13822_), .B(_13815_), .C(_13820_), .Y(_13832_) );
	NAND3X1 NAND3X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_13832_), .B(_13829_), .C(_13831_), .Y(_13833_) );
	NAND3X1 NAND3X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_13828_), .B(_13833_), .C(_13792_), .Y(_13834_) );
	NOR3X1 NOR3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_13520_), .B(_13510_), .C(_13516_), .Y(_13835_) );
	AOI21X1 AOI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .B(_13530_), .C(_13835_), .Y(_13836_) );
	AOI22X1 AOI22X1_320 ( .gnd(gnd), .vdd(vdd), .A(_13799_), .B(_13803_), .C(_13832_), .D(_13831_), .Y(_13837_) );
	AOI21X1 AOI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_13827_), .B(_13821_), .C(_13804_), .Y(_13838_) );
	OAI21X1 OAI21X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_13837_), .B(_13838_), .C(_13836_), .Y(_13839_) );
	NAND3X1 NAND3X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_13834_), .B(_13790_), .C(_13839_), .Y(_13840_) );
	NAND3X1 NAND3X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_13765_), .B(_13787_), .C(_13788_), .Y(_13842_) );
	OAI21X1 OAI21X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_13780_), .B(_13783_), .C(_13785_), .Y(_13843_) );
	NAND2X1 NAND2X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_13842_), .B(_13843_), .Y(_13844_) );
	OAI21X1 OAI21X1_2978 ( .gnd(gnd), .vdd(vdd), .A(_13837_), .B(_13838_), .C(_13792_), .Y(_13845_) );
	NAND3X1 NAND3X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_13828_), .B(_13833_), .C(_13836_), .Y(_13846_) );
	NAND3X1 NAND3X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_13844_), .B(_13846_), .C(_13845_), .Y(_13847_) );
	NAND3X1 NAND3X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_13840_), .B(_13762_), .C(_13847_), .Y(_13848_) );
	NOR3X1 NOR3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13531_), .C(_13534_), .Y(_13849_) );
	AOI21X1 AOI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_13544_), .B(_13547_), .C(_13849_), .Y(_13850_) );
	AOI22X1 AOI22X1_321 ( .gnd(gnd), .vdd(vdd), .A(_13784_), .B(_13789_), .C(_13846_), .D(_13845_), .Y(_13851_) );
	AOI22X1 AOI22X1_322 ( .gnd(gnd), .vdd(vdd), .A(_13842_), .B(_13843_), .C(_13834_), .D(_13839_), .Y(_13853_) );
	OAI21X1 OAI21X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_13851_), .B(_13853_), .C(_13850_), .Y(_13854_) );
	NAND3X1 NAND3X1_2958 ( .gnd(gnd), .vdd(vdd), .A(_13848_), .B(_13854_), .C(_13760_), .Y(_13855_) );
	NAND3X1 NAND3X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_13709_), .B(_13757_), .C(_13758_), .Y(_13856_) );
	OAI21X1 OAI21X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_13749_), .B(_13754_), .C(_13756_), .Y(_13857_) );
	NAND2X1 NAND2X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_13856_), .B(_13857_), .Y(_13858_) );
	OAI21X1 OAI21X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_13851_), .B(_13853_), .C(_13762_), .Y(_13859_) );
	NAND3X1 NAND3X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_13840_), .B(_13847_), .C(_13850_), .Y(_13860_) );
	NAND3X1 NAND3X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_13859_), .B(_13860_), .C(_13858_), .Y(_13861_) );
	NAND3X1 NAND3X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_13855_), .B(_13861_), .C(_13708_), .Y(_13862_) );
	AOI21X1 AOI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_13564_), .B(_13560_), .C(_13567_), .Y(_13864_) );
	AOI22X1 AOI22X1_323 ( .gnd(gnd), .vdd(vdd), .A(_13755_), .B(_13759_), .C(_13859_), .D(_13860_), .Y(_13865_) );
	AOI22X1 AOI22X1_324 ( .gnd(gnd), .vdd(vdd), .A(_13856_), .B(_13857_), .C(_13848_), .D(_13854_), .Y(_13866_) );
	OAI21X1 OAI21X1_2982 ( .gnd(gnd), .vdd(vdd), .A(_13866_), .B(_13865_), .C(_13864_), .Y(_13867_) );
	NAND3X1 NAND3X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_13862_), .B(_13867_), .C(_13707_), .Y(_13868_) );
	NAND3X1 NAND3X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_13703_), .B(_13696_), .C(_13701_), .Y(_13869_) );
	NAND3X1 NAND3X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_13625_), .B(_13704_), .C(_13705_), .Y(_13870_) );
	NAND2X1 NAND2X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_13869_), .B(_13870_), .Y(_13871_) );
	OAI21X1 OAI21X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_13866_), .B(_13865_), .C(_13708_), .Y(_13872_) );
	NAND3X1 NAND3X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_13855_), .B(_13861_), .C(_13864_), .Y(_13873_) );
	NAND3X1 NAND3X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_13872_), .B(_13873_), .C(_13871_), .Y(_13875_) );
	NAND3X1 NAND3X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_13868_), .B(_13875_), .C(_13624_), .Y(_13876_) );
	AOI21X1 AOI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_13575_), .B(_13577_), .C(_13584_), .Y(_13877_) );
	AOI21X1 AOI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_13873_), .B(_13872_), .C(_13871_), .Y(_13878_) );
	AOI21X1 AOI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_13862_), .C(_13707_), .Y(_13879_) );
	OAI21X1 OAI21X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_13879_), .B(_13878_), .C(_13877_), .Y(_13880_) );
	NAND3X1 NAND3X1_2969 ( .gnd(gnd), .vdd(vdd), .A(_13623_), .B(_13880_), .C(_13876_), .Y(_13881_) );
	INVX1 INVX1_1887 ( .gnd(gnd), .vdd(vdd), .A(_13623_), .Y(_13882_) );
	NOR3X1 NOR3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_13879_), .B(_13878_), .C(_13877_), .Y(_13883_) );
	AOI21X1 AOI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_13868_), .B(_13875_), .C(_13624_), .Y(_13884_) );
	OAI21X1 OAI21X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_13884_), .B(_13883_), .C(_13882_), .Y(_13886_) );
	NAND3X1 NAND3X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .B(_13886_), .C(_13615_), .Y(_13887_) );
	INVX1 INVX1_1888 ( .gnd(gnd), .vdd(vdd), .A(_13590_), .Y(_13888_) );
	AOI21X1 AOI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_13589_), .B(_13591_), .C(_13888_), .Y(_13889_) );
	INVX1 INVX1_1889 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .Y(_13890_) );
	AOI21X1 AOI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_13876_), .B(_13880_), .C(_13623_), .Y(_13891_) );
	OAI21X1 OAI21X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_13891_), .B(_13890_), .C(_13889_), .Y(_13892_) );
	NAND3X1 NAND3X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_13892_), .B(_13887_), .C(_13614_), .Y(_13893_) );
	OAI21X1 OAI21X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_13891_), .B(_13890_), .C(_13615_), .Y(_13894_) );
	NAND3X1 NAND3X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .B(_13886_), .C(_13889_), .Y(_13895_) );
	NAND3X1 NAND3X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_13603_), .B(_13895_), .C(_13894_), .Y(_13897_) );
	NAND3X1 NAND3X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_13897_), .B(_13893_), .C(_13613_), .Y(_13898_) );
	AOI21X1 AOI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_13894_), .B(_13895_), .C(_13603_), .Y(_13899_) );
	AOI21X1 AOI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_13887_), .B(_13892_), .C(_13614_), .Y(_13900_) );
	OAI21X1 OAI21X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_13899_), .B(_13900_), .C(_13607_), .Y(_13901_) );
	NAND2X1 NAND2X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_13901_), .B(_13898_), .Y(_13902_) );
	XNOR2X1 XNOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_13612_), .B(_13902_), .Y(mulOut_21_) );
	OAI21X1 OAI21X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_13899_), .B(_13900_), .C(_13613_), .Y(_13903_) );
	NAND2X1 NAND2X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_13897_), .B(_13893_), .Y(_13904_) );
	OAI21X1 OAI21X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_13613_), .B(_13904_), .C(_13606_), .Y(_13905_) );
	NAND2X1 NAND2X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_13903_), .B(_13905_), .Y(_13907_) );
	OAI21X1 OAI21X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .B(_12311_), .C(_12307_), .Y(_13908_) );
	OAI21X1 OAI21X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12305_), .C(_12312_), .Y(_13909_) );
	NAND3X1 NAND3X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_12327_), .B(_13909_), .C(_13908_), .Y(_13910_) );
	OAI21X1 OAI21X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12305_), .C(_12328_), .Y(_13911_) );
	NAND2X1 NAND2X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_13911_), .B(_13910_), .Y(_13912_) );
	AOI21X1 AOI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_11937_), .B(_12315_), .C(_13912_), .Y(_13913_) );
	NOR2X1 NOR2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_17309_), .B(_17310_), .Y(_13914_) );
	NAND3X1 NAND3X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12315_), .C(_13914_), .Y(_13915_) );
	AOI21X1 AOI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_13915_), .B(_13913_), .C(_13321_), .Y(_13916_) );
	AOI21X1 AOI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_12785_), .B(_12784_), .C(_12543_), .Y(_13918_) );
	AOI21X1 AOI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_12556_), .B(_12789_), .C(_13918_), .Y(_13919_) );
	AOI21X1 AOI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_13051_), .B(_13050_), .C(_13049_), .Y(_13920_) );
	AOI21X1 AOI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_13044_), .B(_13047_), .C(_12777_), .Y(_13921_) );
	OAI22X1 OAI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(_13920_), .B(_13921_), .C(_13315_), .D(_13312_), .Y(_13922_) );
	NAND2X1 NAND2X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_13322_), .B(_13324_), .Y(_13923_) );
	OAI21X1 OAI21X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_13919_), .B(_13922_), .C(_13923_), .Y(_13924_) );
	AOI21X1 AOI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_13898_), .B(_13901_), .C(_13610_), .Y(_13925_) );
	OAI21X1 OAI21X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_13924_), .B(_13916_), .C(_13925_), .Y(_13926_) );
	NAND2X1 NAND2X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_13907_), .B(_13926_), .Y(_13927_) );
	NAND2X1 NAND2X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_13881_), .B(_13886_), .Y(_13929_) );
	NOR2X1 NOR2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_13889_), .B(_13929_), .Y(_13930_) );
	OAI21X1 OAI21X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_13882_), .B(_13884_), .C(_13876_), .Y(_13931_) );
	OAI21X1 OAI21X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13639_), .C(_13650_), .Y(_13932_) );
	INVX1 INVX1_1890 ( .gnd(gnd), .vdd(vdd), .A(_13932_), .Y(_13933_) );
	NAND2X1 NAND2X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_13696_), .B(_13869_), .Y(_13934_) );
	OR2X2 OR2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_13934_), .B(_13933_), .Y(_13935_) );
	NAND2X1 NAND2X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_13933_), .B(_13934_), .Y(_13936_) );
	NAND2X1 NAND2X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_13936_), .B(_13935_), .Y(_13937_) );
	AOI21X1 AOI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_13855_), .B(_13861_), .C(_13708_), .Y(_13938_) );
	OAI21X1 OAI21X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_13938_), .B(_13871_), .C(_13862_), .Y(_13940_) );
	INVX1 INVX1_1891 ( .gnd(gnd), .vdd(vdd), .A(_13681_), .Y(_13941_) );
	NOR2X1 NOR2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_13941_), .B(_13697_), .Y(_13942_) );
	AOI22X1 AOI22X1_325 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf3), .B(adder_bOperand_22_bF_buf3), .C(aOperand_frameOut_1_bF_buf2), .D(adder_bOperand_21_bF_buf2), .Y(_13943_) );
	NAND2X1 NAND2X1_2808 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf1), .B(adder_bOperand_22_bF_buf2), .Y(_13944_) );
	NOR2X1 NOR2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13944_), .Y(_13945_) );
	AOI22X1 AOI22X1_326 ( .gnd(gnd), .vdd(vdd), .A(_13641_), .B(_13642_), .C(_13631_), .D(_13635_), .Y(_13946_) );
	INVX1 INVX1_1892 ( .gnd(gnd), .vdd(vdd), .A(_13946_), .Y(_13947_) );
	NOR2X1 NOR2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf3), .B(_13334_), .Y(_13948_) );
	NAND2X1 NAND2X1_2809 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf0), .B(adder_bOperand_18_bF_buf3), .Y(_13949_) );
	NOR2X1 NOR2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_13634_), .B(_13949_), .Y(_13951_) );
	INVX1 INVX1_1893 ( .gnd(gnd), .vdd(vdd), .A(_13951_), .Y(_13952_) );
	OAI21X1 OAI21X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf1), .B(_13338_), .C(_13634_), .Y(_13953_) );
	NAND3X1 NAND3X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_13948_), .B(_13953_), .C(_13952_), .Y(_13954_) );
	NAND3X1 NAND3X1_2978 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf4), .B(adder_bOperand_18_bF_buf2), .C(_13634_), .Y(_13955_) );
	NAND3X1 NAND3X1_2979 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf3), .B(adder_bOperand_19_bF_buf2), .C(_13949_), .Y(_13956_) );
	AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_13955_), .B(_13956_), .Y(_13957_) );
	OAI21X1 OAI21X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf2), .B(_13334_), .C(_13957_), .Y(_13958_) );
	AOI21X1 AOI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_13958_), .B(_13954_), .C(_13947_), .Y(_13959_) );
	INVX1 INVX1_1894 ( .gnd(gnd), .vdd(vdd), .A(_13948_), .Y(_13960_) );
	AOI21X1 AOI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_13955_), .B(_13956_), .C(_13960_), .Y(_13962_) );
	AOI21X1 AOI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_13952_), .B(_13953_), .C(_13948_), .Y(_13963_) );
	NOR3X1 NOR3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_13946_), .B(_13962_), .C(_13963_), .Y(_13964_) );
	OAI22X1 OAI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(_13943_), .B(_13945_), .C(_13959_), .D(_13964_), .Y(_13965_) );
	NOR2X1 NOR2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_13943_), .B(_13945_), .Y(_13966_) );
	OAI21X1 OAI21X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_13962_), .B(_13963_), .C(_13946_), .Y(_13967_) );
	NAND3X1 NAND3X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_13947_), .B(_13954_), .C(_13958_), .Y(_13968_) );
	NAND3X1 NAND3X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_13966_), .B(_13968_), .C(_13967_), .Y(_13969_) );
	AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_13969_), .Y(_13970_) );
	OAI21X1 OAI21X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_13675_), .B(_13679_), .C(_13670_), .Y(_13971_) );
	OAI21X1 OAI21X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .B(_13665_), .C(_13660_), .Y(_13973_) );
	NAND2X1 NAND2X1_2810 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf3), .B(adder_bOperand_17_bF_buf0), .Y(_13974_) );
	INVX1 INVX1_1895 ( .gnd(gnd), .vdd(vdd), .A(_13974_), .Y(_13975_) );
	AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf0), .B(adder_bOperand_15_bF_buf4), .Y(_13976_) );
	NAND2X1 NAND2X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_13659_), .B(_13976_), .Y(_13977_) );
	NAND2X1 NAND2X1_2812 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf4), .B(adder_bOperand_15_bF_buf3), .Y(_13978_) );
	OAI21X1 OAI21X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf1), .B(_12342_), .C(_13978_), .Y(_13979_) );
	NAND3X1 NAND3X1_2982 ( .gnd(gnd), .vdd(vdd), .A(_13975_), .B(_13979_), .C(_13977_), .Y(_13980_) );
	NAND2X1 NAND2X1_2813 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf3), .B(adder_bOperand_16_bF_buf0), .Y(_13981_) );
	NOR2X1 NOR2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_13663_), .B(_13981_), .Y(_13982_) );
	NOR2X1 NOR2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_13659_), .B(_13976_), .Y(_13984_) );
	OAI21X1 OAI21X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_13982_), .B(_13984_), .C(_13974_), .Y(_13985_) );
	AOI21X1 AOI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_13715_), .B(_13711_), .C(_13713_), .Y(_13986_) );
	INVX1 INVX1_1896 ( .gnd(gnd), .vdd(vdd), .A(_13986_), .Y(_13987_) );
	NAND3X1 NAND3X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .B(_13985_), .C(_13987_), .Y(_13988_) );
	INVX1 INVX1_1897 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .Y(_13989_) );
	AOI21X1 AOI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_13977_), .B(_13979_), .C(_13975_), .Y(_13990_) );
	OAI21X1 OAI21X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_13990_), .B(_13989_), .C(_13986_), .Y(_13991_) );
	NAND3X1 NAND3X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_13973_), .B(_13988_), .C(_13991_), .Y(_13992_) );
	INVX1 INVX1_1898 ( .gnd(gnd), .vdd(vdd), .A(_13973_), .Y(_13993_) );
	NAND2X1 NAND2X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .B(_13985_), .Y(_13995_) );
	NOR2X1 NOR2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_13986_), .B(_13995_), .Y(_13996_) );
	AOI21X1 AOI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_13985_), .B(_13980_), .C(_13987_), .Y(_13997_) );
	OAI21X1 OAI21X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_13997_), .B(_13996_), .C(_13993_), .Y(_13998_) );
	NAND3X1 NAND3X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_13992_), .B(_13971_), .C(_13998_), .Y(_13999_) );
	AOI21X1 AOI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_13673_), .B(_13656_), .C(_13678_), .Y(_14000_) );
	NAND3X1 NAND3X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .B(_13986_), .C(_13985_), .Y(_14001_) );
	OAI21X1 OAI21X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_13990_), .B(_13989_), .C(_13987_), .Y(_14002_) );
	AOI21X1 AOI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_14002_), .B(_14001_), .C(_13993_), .Y(_14003_) );
	AOI21X1 AOI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_13991_), .B(_13988_), .C(_13973_), .Y(_14004_) );
	OAI21X1 OAI21X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_14003_), .B(_14004_), .C(_14000_), .Y(_14006_) );
	NAND3X1 NAND3X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_14006_), .B(_13999_), .C(_13970_), .Y(_14007_) );
	NAND2X1 NAND2X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_13969_), .B(_13965_), .Y(_14008_) );
	OAI21X1 OAI21X1_3010 ( .gnd(gnd), .vdd(vdd), .A(_14003_), .B(_14004_), .C(_13971_), .Y(_14009_) );
	NAND3X1 NAND3X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_14000_), .B(_13992_), .C(_13998_), .Y(_14010_) );
	NAND3X1 NAND3X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_14008_), .B(_14009_), .C(_14010_), .Y(_14011_) );
	OAI21X1 OAI21X1_3011 ( .gnd(gnd), .vdd(vdd), .A(_13749_), .B(_13756_), .C(_13758_), .Y(_14012_) );
	NAND3X1 NAND3X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_14011_), .B(_14012_), .C(_14007_), .Y(_14013_) );
	AOI21X1 AOI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_14010_), .B(_14009_), .C(_14008_), .Y(_14014_) );
	AOI22X1 AOI22X1_327 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_13969_), .C(_14006_), .D(_13999_), .Y(_14015_) );
	AOI21X1 AOI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_13709_), .B(_13757_), .C(_13754_), .Y(_14017_) );
	OAI21X1 OAI21X1_3012 ( .gnd(gnd), .vdd(vdd), .A(_14015_), .B(_14014_), .C(_14017_), .Y(_14018_) );
	NAND3X1 NAND3X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_13942_), .B(_14013_), .C(_14018_), .Y(_14019_) );
	NAND2X1 NAND2X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_13681_), .B(_13690_), .Y(_14020_) );
	NAND3X1 NAND3X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_14017_), .B(_14011_), .C(_14007_), .Y(_14021_) );
	OAI21X1 OAI21X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_14015_), .B(_14014_), .C(_14012_), .Y(_14022_) );
	NAND3X1 NAND3X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_14020_), .B(_14021_), .C(_14022_), .Y(_14023_) );
	NAND2X1 NAND2X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_14019_), .B(_14023_), .Y(_14024_) );
	AOI21X1 AOI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_13847_), .B(_13840_), .C(_13762_), .Y(_14025_) );
	OAI21X1 OAI21X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_14025_), .B(_13858_), .C(_13848_), .Y(_14026_) );
	AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_13743_), .B(_13735_), .Y(_14027_) );
	NOR2X1 NOR2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_12365_), .Y(_14028_) );
	NAND2X1 NAND2X1_2818 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf4), .B(adder_bOperand_13_bF_buf0), .Y(_14029_) );
	NAND2X1 NAND2X1_2819 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf2), .B(adder_bOperand_13_bF_buf3), .Y(_14030_) );
	OAI21X1 OAI21X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_17157_), .C(_14030_), .Y(_14031_) );
	OAI21X1 OAI21X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_13712_), .B(_14029_), .C(_14031_), .Y(_14032_) );
	XNOR2X1 XNOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_14032_), .B(_14028_), .Y(_14033_) );
	AOI21X1 AOI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_13729_), .B(_13724_), .C(_13732_), .Y(_14034_) );
	INVX1 INVX1_1899 ( .gnd(gnd), .vdd(vdd), .A(_14034_), .Y(_14035_) );
	NOR2X1 NOR2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_17022__bF_buf3), .Y(_14036_) );
	NAND2X1 NAND2X1_2820 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf3), .B(aOperand_frameOut_13_bF_buf4), .Y(_14038_) );
	INVX1 INVX1_1900 ( .gnd(gnd), .vdd(vdd), .A(_14038_), .Y(_14039_) );
	NAND2X1 NAND2X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_13726_), .B(_14039_), .Y(_14040_) );
	NAND2X1 NAND2X1_2822 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf0), .B(aOperand_frameOut_13_bF_buf3), .Y(_14041_) );
	OAI21X1 OAI21X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_16887_), .B(_17236__bF_buf3), .C(_14041_), .Y(_14042_) );
	NAND3X1 NAND3X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_14036_), .B(_14042_), .C(_14040_), .Y(_14043_) );
	OAI21X1 OAI21X1_3018 ( .gnd(gnd), .vdd(vdd), .A(_13731_), .B(_14038_), .C(_14042_), .Y(_14044_) );
	OAI21X1 OAI21X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_17022__bF_buf2), .C(_14044_), .Y(_14045_) );
	NAND3X1 NAND3X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_14043_), .B(_14045_), .C(_14035_), .Y(_14046_) );
	INVX1 INVX1_1901 ( .gnd(gnd), .vdd(vdd), .A(_14036_), .Y(_14047_) );
	NOR2X1 NOR2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_14047_), .B(_14044_), .Y(_14050_) );
	AOI21X1 AOI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_14040_), .B(_14042_), .C(_14036_), .Y(_14051_) );
	OAI21X1 OAI21X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_14051_), .B(_14050_), .C(_14034_), .Y(_14052_) );
	NAND3X1 NAND3X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_14033_), .B(_14046_), .C(_14052_), .Y(_14053_) );
	INVX1 INVX1_1902 ( .gnd(gnd), .vdd(vdd), .A(_14028_), .Y(_14054_) );
	OR2X2 OR2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_14032_), .B(_14054_), .Y(_14055_) );
	OAI21X1 OAI21X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_12365_), .C(_14032_), .Y(_14056_) );
	NAND2X1 NAND2X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_14056_), .B(_14055_), .Y(_14057_) );
	OAI21X1 OAI21X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_14051_), .B(_14050_), .C(_14035_), .Y(_14058_) );
	NAND3X1 NAND3X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_14034_), .B(_14043_), .C(_14045_), .Y(_14059_) );
	NAND3X1 NAND3X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_14059_), .B(_14057_), .C(_14058_), .Y(_14061_) );
	OAI21X1 OAI21X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_13780_), .B(_13785_), .C(_13788_), .Y(_14062_) );
	NAND3X1 NAND3X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_14062_), .B(_14053_), .C(_14061_), .Y(_14063_) );
	AOI21X1 AOI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_14058_), .B(_14059_), .C(_14057_), .Y(_14064_) );
	AOI21X1 AOI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_14052_), .B(_14046_), .C(_14033_), .Y(_14065_) );
	AOI21X1 AOI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_13787_), .B(_13765_), .C(_13783_), .Y(_14066_) );
	OAI21X1 OAI21X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_14065_), .B(_14064_), .C(_14066_), .Y(_14067_) );
	NAND3X1 NAND3X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_14027_), .B(_14063_), .C(_14067_), .Y(_14068_) );
	NAND2X1 NAND2X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_13735_), .B(_13743_), .Y(_14069_) );
	NAND3X1 NAND3X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_14066_), .B(_14053_), .C(_14061_), .Y(_14070_) );
	OAI21X1 OAI21X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_14065_), .B(_14064_), .C(_14062_), .Y(_14072_) );
	NAND3X1 NAND3X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_14069_), .B(_14070_), .C(_14072_), .Y(_14073_) );
	NAND2X1 NAND2X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_14068_), .B(_14073_), .Y(_14074_) );
	AOI21X1 AOI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_13833_), .B(_13828_), .C(_13792_), .Y(_14075_) );
	OAI21X1 OAI21X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_14075_), .B(_13844_), .C(_13834_), .Y(_14076_) );
	NAND2X1 NAND2X1_2826 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf2), .B(aOperand_frameOut_15_bF_buf3), .Y(_14077_) );
	OAI21X1 OAI21X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .B(_14077_), .C(_13771_), .Y(_14078_) );
	INVX1 INVX1_1903 ( .gnd(gnd), .vdd(vdd), .A(_14078_), .Y(_14079_) );
	NAND2X1 NAND2X1_2827 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf3), .B(aOperand_frameOut_14_bF_buf2), .Y(_14080_) );
	INVX1 INVX1_1904 ( .gnd(gnd), .vdd(vdd), .A(_14080_), .Y(_14081_) );
	AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf2), .B(aOperand_frameOut_16_bF_buf4), .Y(_14083_) );
	NAND2X1 NAND2X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_13768_), .B(_14083_), .Y(_14084_) );
	OAI21X1 OAI21X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf1), .B(_12461_), .C(_14077_), .Y(_14085_) );
	NAND3X1 NAND3X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_14081_), .B(_14085_), .C(_14084_), .Y(_14086_) );
	OAI21X1 OAI21X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_13830_), .B(_12233_), .C(_14083_), .Y(_14087_) );
	OAI21X1 OAI21X1_3030 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf0), .B(_12461_), .C(_13768_), .Y(_14088_) );
	NAND3X1 NAND3X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_14080_), .B(_14087_), .C(_14088_), .Y(_14089_) );
	NOR2X1 NOR2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_13777_), .B(_13794_), .Y(_14090_) );
	OAI21X1 OAI21X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_13793_), .B(_14090_), .C(_13795_), .Y(_14091_) );
	NAND3X1 NAND3X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_14086_), .B(_14089_), .C(_14091_), .Y(_14092_) );
	AOI21X1 AOI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_14087_), .B(_14088_), .C(_14080_), .Y(_14094_) );
	AOI21X1 AOI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_14084_), .B(_14085_), .C(_14081_), .Y(_14095_) );
	NAND2X1 NAND2X1_2829 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf5), .B(aOperand_frameOut_18_bF_buf4), .Y(_14096_) );
	INVX1 INVX1_1905 ( .gnd(gnd), .vdd(vdd), .A(_14096_), .Y(_14097_) );
	AOI22X1 AOI22X1_328 ( .gnd(gnd), .vdd(vdd), .A(_13492_), .B(_14097_), .C(_13800_), .D(_13798_), .Y(_14098_) );
	OAI21X1 OAI21X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_14095_), .B(_14094_), .C(_14098_), .Y(_14099_) );
	NAND3X1 NAND3X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_14092_), .B(_14099_), .C(_14079_), .Y(_14100_) );
	NAND3X1 NAND3X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_14086_), .B(_14098_), .C(_14089_), .Y(_14101_) );
	OAI21X1 OAI21X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_14095_), .B(_14094_), .C(_14091_), .Y(_14102_) );
	NAND3X1 NAND3X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_14078_), .B(_14101_), .C(_14102_), .Y(_14103_) );
	NAND2X1 NAND2X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_14103_), .B(_14100_), .Y(_14105_) );
	AOI21X1 AOI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_13820_), .B(_13815_), .C(_13806_), .Y(_14106_) );
	OAI21X1 OAI21X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_13829_), .B(_14106_), .C(_13821_), .Y(_14107_) );
	NOR2X1 NOR2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf3), .B(_12708_), .Y(_14108_) );
	INVX1 INVX1_1906 ( .gnd(gnd), .vdd(vdd), .A(_14108_), .Y(_14109_) );
	NAND2X1 NAND2X1_2831 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf5), .B(aOperand_frameOut_19_bF_buf0), .Y(_14110_) );
	NOR2X1 NOR2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_14096_), .B(_14110_), .Y(_14111_) );
	INVX1 INVX1_1907 ( .gnd(gnd), .vdd(vdd), .A(_14111_), .Y(_14112_) );
	OAI21X1 OAI21X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf0), .B(_13224_), .C(_14096_), .Y(_14113_) );
	NAND3X1 NAND3X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_14109_), .B(_14113_), .C(_14112_), .Y(_14114_) );
	AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_14096_), .B(_14110_), .Y(_14116_) );
	OAI21X1 OAI21X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_14111_), .B(_14116_), .C(_14108_), .Y(_14117_) );
	NAND2X1 NAND2X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_14117_), .B(_14114_), .Y(_14118_) );
	OAI21X1 OAI21X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_13807_), .B(_13818_), .C(_13811_), .Y(_14119_) );
	NAND2X1 NAND2X1_2833 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf5), .B(aOperand_frameOut_20_bF_buf4), .Y(_14120_) );
	INVX1 INVX1_1908 ( .gnd(gnd), .vdd(vdd), .A(_14120_), .Y(_14121_) );
	AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf1), .B(aOperand_frameOut_21_bF_buf0), .Y(_14122_) );
	AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .B(aOperand_frameOut_22_bF_buf0), .Y(_14123_) );
	NAND2X1 NAND2X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_14122_), .B(_14123_), .Y(_14124_) );
	INVX4 INVX4_23 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_22_bF_buf3), .Y(_14125_) );
	NAND2X1 NAND2X1_2835 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf0), .B(aOperand_frameOut_21_bF_buf4), .Y(_14127_) );
	OAI21X1 OAI21X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf0), .B(_14125_), .C(_14127_), .Y(_14128_) );
	NAND3X1 NAND3X1_3010 ( .gnd(gnd), .vdd(vdd), .A(_14121_), .B(_14128_), .C(_14124_), .Y(_14129_) );
	NAND3X1 NAND3X1_3011 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_22_bF_buf2), .C(_14127_), .Y(_14130_) );
	NAND2X1 NAND2X1_2836 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_22_bF_buf1), .Y(_14131_) );
	NAND3X1 NAND3X1_3012 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf6), .B(aOperand_frameOut_21_bF_buf3), .C(_14131_), .Y(_14132_) );
	NAND3X1 NAND3X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_14120_), .B(_14130_), .C(_14132_), .Y(_14133_) );
	NAND3X1 NAND3X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_14129_), .B(_14133_), .C(_14119_), .Y(_14134_) );
	AOI21X1 AOI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_13814_), .B(_13809_), .C(_13817_), .Y(_14135_) );
	AOI21X1 AOI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_14130_), .B(_14132_), .C(_14120_), .Y(_14136_) );
	AOI22X1 AOI22X1_329 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .B(aOperand_frameOut_20_bF_buf3), .C(_14128_), .D(_14124_), .Y(_14138_) );
	OAI21X1 OAI21X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_14136_), .B(_14138_), .C(_14135_), .Y(_14139_) );
	NAND3X1 NAND3X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_14134_), .B(_14139_), .C(_14118_), .Y(_14140_) );
	NAND3X1 NAND3X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_14108_), .B(_14113_), .C(_14112_), .Y(_14141_) );
	OAI21X1 OAI21X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_14111_), .B(_14116_), .C(_14109_), .Y(_14142_) );
	NAND2X1 NAND2X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_14142_), .B(_14141_), .Y(_14143_) );
	OAI21X1 OAI21X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_14136_), .B(_14138_), .C(_14119_), .Y(_14144_) );
	NAND3X1 NAND3X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_14133_), .B(_14129_), .C(_14135_), .Y(_14145_) );
	NAND3X1 NAND3X1_3018 ( .gnd(gnd), .vdd(vdd), .A(_14145_), .B(_14144_), .C(_14143_), .Y(_14146_) );
	NAND3X1 NAND3X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_14140_), .B(_14146_), .C(_14107_), .Y(_14147_) );
	NOR3X1 NOR3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_13822_), .B(_13825_), .C(_13826_), .Y(_14149_) );
	AOI21X1 AOI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_13804_), .B(_13827_), .C(_14149_), .Y(_14150_) );
	AOI21X1 AOI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_14144_), .B(_14145_), .C(_14143_), .Y(_14151_) );
	AOI21X1 AOI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_14139_), .B(_14134_), .C(_14118_), .Y(_14152_) );
	OAI21X1 OAI21X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_14151_), .B(_14152_), .C(_14150_), .Y(_14153_) );
	NAND3X1 NAND3X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_14105_), .B(_14147_), .C(_14153_), .Y(_14154_) );
	NAND3X1 NAND3X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_14078_), .B(_14092_), .C(_14099_), .Y(_14155_) );
	NAND3X1 NAND3X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_14101_), .B(_14102_), .C(_14079_), .Y(_14156_) );
	NAND2X1 NAND2X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_14155_), .B(_14156_), .Y(_14157_) );
	OAI21X1 OAI21X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_14151_), .B(_14152_), .C(_14107_), .Y(_14158_) );
	NAND3X1 NAND3X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_14140_), .B(_14146_), .C(_14150_), .Y(_14160_) );
	NAND3X1 NAND3X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_14157_), .B(_14160_), .C(_14158_), .Y(_14161_) );
	NAND3X1 NAND3X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_14154_), .B(_14076_), .C(_14161_), .Y(_14162_) );
	INVX1 INVX1_1909 ( .gnd(gnd), .vdd(vdd), .A(_13834_), .Y(_14163_) );
	AOI21X1 AOI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_13790_), .B(_13839_), .C(_14163_), .Y(_14164_) );
	AOI22X1 AOI22X1_330 ( .gnd(gnd), .vdd(vdd), .A(_14100_), .B(_14103_), .C(_14160_), .D(_14158_), .Y(_14165_) );
	AOI22X1 AOI22X1_331 ( .gnd(gnd), .vdd(vdd), .A(_14155_), .B(_14156_), .C(_14147_), .D(_14153_), .Y(_14166_) );
	OAI21X1 OAI21X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_14165_), .B(_14166_), .C(_14164_), .Y(_14167_) );
	NAND3X1 NAND3X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_14162_), .B(_14167_), .C(_14074_), .Y(_14168_) );
	NAND3X1 NAND3X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_14069_), .B(_14063_), .C(_14067_), .Y(_14169_) );
	NAND3X1 NAND3X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_14027_), .B(_14070_), .C(_14072_), .Y(_14171_) );
	NAND2X1 NAND2X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_14169_), .B(_14171_), .Y(_14172_) );
	OAI21X1 OAI21X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_14165_), .B(_14166_), .C(_14076_), .Y(_14173_) );
	NAND3X1 NAND3X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_14154_), .B(_14161_), .C(_14164_), .Y(_14174_) );
	NAND3X1 NAND3X1_3030 ( .gnd(gnd), .vdd(vdd), .A(_14173_), .B(_14174_), .C(_14172_), .Y(_14175_) );
	NAND3X1 NAND3X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_14168_), .B(_14175_), .C(_14026_), .Y(_14176_) );
	INVX1 INVX1_1910 ( .gnd(gnd), .vdd(vdd), .A(_13848_), .Y(_14177_) );
	AOI21X1 AOI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_13760_), .B(_13854_), .C(_14177_), .Y(_14178_) );
	AOI22X1 AOI22X1_332 ( .gnd(gnd), .vdd(vdd), .A(_14068_), .B(_14073_), .C(_14173_), .D(_14174_), .Y(_14179_) );
	AOI22X1 AOI22X1_333 ( .gnd(gnd), .vdd(vdd), .A(_14169_), .B(_14171_), .C(_14162_), .D(_14167_), .Y(_14180_) );
	OAI21X1 OAI21X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_14180_), .B(_14179_), .C(_14178_), .Y(_14182_) );
	NAND3X1 NAND3X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_14176_), .B(_14182_), .C(_14024_), .Y(_14183_) );
	NAND3X1 NAND3X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_14020_), .B(_14013_), .C(_14018_), .Y(_14184_) );
	NAND3X1 NAND3X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_13942_), .B(_14021_), .C(_14022_), .Y(_14185_) );
	NAND2X1 NAND2X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_14185_), .B(_14184_), .Y(_14186_) );
	OAI21X1 OAI21X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_14180_), .B(_14179_), .C(_14026_), .Y(_14187_) );
	NAND3X1 NAND3X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_14168_), .B(_14175_), .C(_14178_), .Y(_14188_) );
	NAND3X1 NAND3X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_14187_), .B(_14188_), .C(_14186_), .Y(_14189_) );
	NAND3X1 NAND3X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_14183_), .B(_14189_), .C(_13940_), .Y(_14190_) );
	NOR3X1 NOR3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_13866_), .B(_13865_), .C(_13864_), .Y(_14191_) );
	AOI21X1 AOI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_13707_), .B(_13867_), .C(_14191_), .Y(_14193_) );
	AOI22X1 AOI22X1_334 ( .gnd(gnd), .vdd(vdd), .A(_14019_), .B(_14023_), .C(_14187_), .D(_14188_), .Y(_14194_) );
	AOI22X1 AOI22X1_335 ( .gnd(gnd), .vdd(vdd), .A(_14184_), .B(_14185_), .C(_14176_), .D(_14182_), .Y(_14195_) );
	OAI21X1 OAI21X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_14195_), .B(_14194_), .C(_14193_), .Y(_14196_) );
	NAND3X1 NAND3X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_13937_), .B(_14190_), .C(_14196_), .Y(_14197_) );
	NAND2X1 NAND2X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_13932_), .B(_13934_), .Y(_14198_) );
	OR2X2 OR2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_13934_), .B(_13932_), .Y(_14199_) );
	NAND2X1 NAND2X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .B(_14199_), .Y(_14200_) );
	OAI21X1 OAI21X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_14195_), .B(_14194_), .C(_13940_), .Y(_14201_) );
	NAND3X1 NAND3X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_14183_), .B(_14189_), .C(_14193_), .Y(_14202_) );
	NAND3X1 NAND3X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_14200_), .B(_14201_), .C(_14202_), .Y(_14204_) );
	NAND3X1 NAND3X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_14197_), .B(_14204_), .C(_13931_), .Y(_14205_) );
	AOI21X1 AOI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_13623_), .B(_13880_), .C(_13883_), .Y(_14206_) );
	AOI21X1 AOI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_14202_), .B(_14201_), .C(_14200_), .Y(_14207_) );
	AOI22X1 AOI22X1_336 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .B(_14199_), .C(_14190_), .D(_14196_), .Y(_14208_) );
	OAI21X1 OAI21X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_14208_), .B(_14207_), .C(_14206_), .Y(_14209_) );
	NAND3X1 NAND3X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_13619_), .B(_14205_), .C(_14209_), .Y(_14210_) );
	OAI21X1 OAI21X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_14208_), .B(_14207_), .C(_13931_), .Y(_14211_) );
	NAND3X1 NAND3X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_14197_), .B(_14204_), .C(_14206_), .Y(_14212_) );
	NAND3X1 NAND3X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .B(_14211_), .C(_14212_), .Y(_14213_) );
	NAND3X1 NAND3X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_14210_), .B(_13930_), .C(_14213_), .Y(_14215_) );
	NAND3X1 NAND3X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .B(_14205_), .C(_14209_), .Y(_14216_) );
	NAND3X1 NAND3X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_13619_), .B(_14211_), .C(_14212_), .Y(_14217_) );
	NAND3X1 NAND3X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_13887_), .B(_14216_), .C(_14217_), .Y(_14218_) );
	NAND3X1 NAND3X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_13893_), .B(_14218_), .C(_14215_), .Y(_14219_) );
	NAND3X1 NAND3X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_13887_), .B(_14210_), .C(_14213_), .Y(_14220_) );
	NAND3X1 NAND3X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_14216_), .B(_13930_), .C(_14217_), .Y(_14221_) );
	NAND3X1 NAND3X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_13899_), .B(_14220_), .C(_14221_), .Y(_14222_) );
	NAND2X1 NAND2X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_14219_), .B(_14222_), .Y(_14223_) );
	AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_13927_), .B(_14223_), .Y(_14224_) );
	NOR2X1 NOR2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_14223_), .B(_13927_), .Y(_14226_) );
	NOR2X1 NOR2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_14226_), .B(_14224_), .Y(mulOut_22_) );
	NAND3X1 NAND3X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_13899_), .B(_14218_), .C(_14215_), .Y(_14227_) );
	INVX1 INVX1_1911 ( .gnd(gnd), .vdd(vdd), .A(_14227_), .Y(_14228_) );
	NOR2X1 NOR2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_14228_), .B(_14224_), .Y(_14229_) );
	AOI21X1 AOI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_14197_), .B(_14204_), .C(_13931_), .Y(_14230_) );
	OAI21X1 OAI21X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .B(_14230_), .C(_14205_), .Y(_14231_) );
	INVX1 INVX1_1912 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .Y(_14232_) );
	AOI21X1 AOI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_14189_), .B(_14183_), .C(_13940_), .Y(_14233_) );
	OAI21X1 OAI21X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_14200_), .B(_14233_), .C(_14190_), .Y(_14234_) );
	NAND2X1 NAND2X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_13968_), .B(_13969_), .Y(_14236_) );
	INVX1 INVX1_1913 ( .gnd(gnd), .vdd(vdd), .A(_14236_), .Y(_14237_) );
	OAI21X1 OAI21X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13944_), .C(_14237_), .Y(_14238_) );
	NAND2X1 NAND2X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_13945_), .B(_13964_), .Y(_14239_) );
	NAND2X1 NAND2X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_14239_), .B(_14238_), .Y(_14240_) );
	NAND2X1 NAND2X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_14013_), .B(_14184_), .Y(_14241_) );
	OR2X2 OR2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_14241_), .B(_14240_), .Y(_14242_) );
	NAND2X1 NAND2X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_14240_), .B(_14241_), .Y(_14243_) );
	NAND2X1 NAND2X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_14243_), .B(_14242_), .Y(_14244_) );
	AOI21X1 AOI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_14175_), .B(_14168_), .C(_14026_), .Y(_14245_) );
	OAI21X1 OAI21X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_14245_), .B(_14186_), .C(_14176_), .Y(_14247_) );
	AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_14007_), .B(_13999_), .Y(_14248_) );
	NAND2X1 NAND2X1_2850 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf2), .B(adder_bOperand_23_), .Y(_14249_) );
	NAND2X1 NAND2X1_2851 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf4), .B(adder_bOperand_21_bF_buf1), .Y(_14250_) );
	XOR2X1 XOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_13944_), .B(_14250_), .Y(_14251_) );
	XNOR2X1 XNOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_14251_), .B(_14249_), .Y(_14252_) );
	INVX1 INVX1_1914 ( .gnd(gnd), .vdd(vdd), .A(_14252_), .Y(_14253_) );
	AOI21X1 AOI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_13953_), .B(_13948_), .C(_13951_), .Y(_14254_) );
	INVX1 INVX1_1915 ( .gnd(gnd), .vdd(vdd), .A(_14254_), .Y(_14255_) );
	NAND2X1 NAND2X1_2852 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .B(adder_bOperand_20_bF_buf3), .Y(_14256_) );
	NAND2X1 NAND2X1_2853 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf2), .B(adder_bOperand_19_bF_buf1), .Y(_14258_) );
	NAND2X1 NAND2X1_2854 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf1), .B(adder_bOperand_18_bF_buf1), .Y(_14259_) );
	OAI21X1 OAI21X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf0), .B(_13067_), .C(_14259_), .Y(_14260_) );
	OAI21X1 OAI21X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_13949_), .B(_14258_), .C(_14260_), .Y(_14261_) );
	OR2X2 OR2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_14261_), .B(_14256_), .Y(_14262_) );
	OAI21X1 OAI21X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_13334_), .C(_14261_), .Y(_14263_) );
	AOI21X1 AOI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_14262_), .B(_14263_), .C(_14255_), .Y(_14264_) );
	NOR2X1 NOR2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_14256_), .B(_14261_), .Y(_14265_) );
	AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_14261_), .B(_14256_), .Y(_14266_) );
	NOR3X1 NOR3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_14254_), .B(_14265_), .C(_14266_), .Y(_14267_) );
	OAI21X1 OAI21X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_14264_), .B(_14267_), .C(_14253_), .Y(_14269_) );
	OAI21X1 OAI21X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_14265_), .B(_14266_), .C(_14254_), .Y(_14270_) );
	NAND3X1 NAND3X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_14255_), .B(_14263_), .C(_14262_), .Y(_14271_) );
	NAND3X1 NAND3X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_14252_), .B(_14271_), .C(_14270_), .Y(_14272_) );
	AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_14269_), .B(_14272_), .Y(_14273_) );
	OAI21X1 OAI21X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_13993_), .B(_13997_), .C(_13988_), .Y(_14274_) );
	OAI21X1 OAI21X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_13974_), .B(_13984_), .C(_13977_), .Y(_14275_) );
	OAI21X1 OAI21X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_12131_), .C(_13981_), .Y(_14276_) );
	NAND2X1 NAND2X1_2855 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf2), .B(adder_bOperand_16_bF_buf3), .Y(_14277_) );
	OAI21X1 OAI21X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_13978_), .B(_14277_), .C(_14276_), .Y(_14278_) );
	OAI21X1 OAI21X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf0), .B(_12566_), .C(_14278_), .Y(_14280_) );
	NOR2X1 NOR2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf3), .B(_12566_), .Y(_14281_) );
	NAND2X1 NAND2X1_2856 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf1), .B(adder_bOperand_15_bF_buf2), .Y(_14282_) );
	OR2X2 OR2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_13981_), .B(_14282_), .Y(_14283_) );
	NAND3X1 NAND3X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_14281_), .B(_14276_), .C(_14283_), .Y(_14284_) );
	INVX1 INVX1_1916 ( .gnd(gnd), .vdd(vdd), .A(_13712_), .Y(_14285_) );
	INVX1 INVX1_1917 ( .gnd(gnd), .vdd(vdd), .A(_14029_), .Y(_14286_) );
	AOI22X1 AOI22X1_337 ( .gnd(gnd), .vdd(vdd), .A(_14285_), .B(_14286_), .C(_14028_), .D(_14031_), .Y(_14287_) );
	INVX1 INVX1_1918 ( .gnd(gnd), .vdd(vdd), .A(_14287_), .Y(_14288_) );
	NAND3X1 NAND3X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_14284_), .B(_14280_), .C(_14288_), .Y(_14289_) );
	AOI21X1 AOI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_14283_), .B(_14276_), .C(_14281_), .Y(_14291_) );
	INVX1 INVX1_1919 ( .gnd(gnd), .vdd(vdd), .A(_14281_), .Y(_14292_) );
	NOR2X1 NOR2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_14292_), .B(_14278_), .Y(_14293_) );
	OAI21X1 OAI21X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_14291_), .B(_14293_), .C(_14287_), .Y(_14294_) );
	NAND3X1 NAND3X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_14275_), .B(_14289_), .C(_14294_), .Y(_14295_) );
	INVX1 INVX1_1920 ( .gnd(gnd), .vdd(vdd), .A(_14275_), .Y(_14296_) );
	NAND3X1 NAND3X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_14284_), .B(_14287_), .C(_14280_), .Y(_14297_) );
	OAI21X1 OAI21X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_14291_), .B(_14293_), .C(_14288_), .Y(_14298_) );
	NAND3X1 NAND3X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_14296_), .B(_14297_), .C(_14298_), .Y(_14299_) );
	NAND3X1 NAND3X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_14295_), .B(_14274_), .C(_14299_), .Y(_14300_) );
	AOI21X1 AOI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_13973_), .B(_13991_), .C(_13996_), .Y(_14302_) );
	AOI21X1 AOI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_14298_), .B(_14297_), .C(_14296_), .Y(_14303_) );
	AOI21X1 AOI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_14294_), .B(_14289_), .C(_14275_), .Y(_14304_) );
	OAI21X1 OAI21X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_14303_), .B(_14304_), .C(_14302_), .Y(_14305_) );
	NAND3X1 NAND3X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_14300_), .B(_14305_), .C(_14273_), .Y(_14306_) );
	NAND2X1 NAND2X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_14272_), .B(_14269_), .Y(_14307_) );
	OAI21X1 OAI21X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_14303_), .B(_14304_), .C(_14274_), .Y(_14308_) );
	NAND3X1 NAND3X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_14295_), .B(_14299_), .C(_14302_), .Y(_14309_) );
	NAND3X1 NAND3X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_14309_), .B(_14308_), .C(_14307_), .Y(_14310_) );
	AOI21X1 AOI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_14061_), .B(_14053_), .C(_14062_), .Y(_14311_) );
	OAI21X1 OAI21X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_14027_), .B(_14311_), .C(_14063_), .Y(_14313_) );
	NAND3X1 NAND3X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_14310_), .B(_14313_), .C(_14306_), .Y(_14314_) );
	AOI21X1 AOI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_14308_), .B(_14309_), .C(_14307_), .Y(_14315_) );
	AOI22X1 AOI22X1_338 ( .gnd(gnd), .vdd(vdd), .A(_14269_), .B(_14272_), .C(_14300_), .D(_14305_), .Y(_14316_) );
	INVX1 INVX1_1921 ( .gnd(gnd), .vdd(vdd), .A(_14063_), .Y(_14317_) );
	AOI21X1 AOI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_14069_), .B(_14067_), .C(_14317_), .Y(_14318_) );
	OAI21X1 OAI21X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_14316_), .B(_14315_), .C(_14318_), .Y(_14319_) );
	NAND3X1 NAND3X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_14314_), .B(_14248_), .C(_14319_), .Y(_14320_) );
	NAND2X1 NAND2X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_13999_), .B(_14007_), .Y(_14321_) );
	NAND3X1 NAND3X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_14310_), .B(_14306_), .C(_14318_), .Y(_14322_) );
	OAI21X1 OAI21X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_14316_), .B(_14315_), .C(_14313_), .Y(_14324_) );
	NAND3X1 NAND3X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .B(_14324_), .C(_14322_), .Y(_14325_) );
	NAND2X1 NAND2X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_14320_), .B(_14325_), .Y(_14326_) );
	AOI21X1 AOI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_14161_), .B(_14154_), .C(_14076_), .Y(_14327_) );
	OAI21X1 OAI21X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_14327_), .B(_14172_), .C(_14162_), .Y(_14328_) );
	AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_14053_), .B(_14046_), .Y(_14329_) );
	NOR2X1 NOR2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf3), .B(_12365_), .Y(_14330_) );
	NOR2X1 NOR2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_17157_), .Y(_14331_) );
	NAND2X1 NAND2X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_14286_), .B(_14331_), .Y(_14332_) );
	OAI21X1 OAI21X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_17157_), .C(_14029_), .Y(_14333_) );
	NAND3X1 NAND3X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_14330_), .B(_14333_), .C(_14332_), .Y(_14335_) );
	NAND2X1 NAND2X1_2861 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf3), .B(adder_bOperand_12_bF_buf2), .Y(_14336_) );
	NAND2X1 NAND2X1_2862 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf1), .B(adder_bOperand_13_bF_buf2), .Y(_14337_) );
	OAI21X1 OAI21X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_14336_), .B(_14337_), .C(_14333_), .Y(_14338_) );
	OAI21X1 OAI21X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf2), .B(_12365_), .C(_14338_), .Y(_14339_) );
	NAND2X1 NAND2X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_14335_), .B(_14339_), .Y(_14340_) );
	INVX1 INVX1_1922 ( .gnd(gnd), .vdd(vdd), .A(_14340_), .Y(_14341_) );
	AOI22X1 AOI22X1_339 ( .gnd(gnd), .vdd(vdd), .A(_14039_), .B(_13726_), .C(_14036_), .D(_14042_), .Y(_14342_) );
	INVX1 INVX1_1923 ( .gnd(gnd), .vdd(vdd), .A(_14342_), .Y(_14343_) );
	NOR2X1 NOR2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf1), .B(_17236__bF_buf2), .Y(_14344_) );
	INVX1 INVX1_1924 ( .gnd(gnd), .vdd(vdd), .A(_14344_), .Y(_14346_) );
	NAND2X1 NAND2X1_2864 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf2), .B(aOperand_frameOut_14_bF_buf1), .Y(_14347_) );
	OAI21X1 OAI21X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf0), .B(_12039_), .C(_14038_), .Y(_14348_) );
	OAI21X1 OAI21X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_14041_), .B(_14347_), .C(_14348_), .Y(_14349_) );
	OR2X2 OR2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_14349_), .B(_14346_), .Y(_14350_) );
	OAI21X1 OAI21X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf0), .B(_17236__bF_buf1), .C(_14349_), .Y(_14351_) );
	NAND3X1 NAND3X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_14351_), .B(_14343_), .C(_14350_), .Y(_14352_) );
	NOR2X1 NOR2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_14346_), .B(_14349_), .Y(_14353_) );
	NAND2X1 NAND2X1_2865 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf4), .B(aOperand_frameOut_14_bF_buf0), .Y(_14354_) );
	INVX1 INVX1_1925 ( .gnd(gnd), .vdd(vdd), .A(_14354_), .Y(_14355_) );
	NAND2X1 NAND2X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_14039_), .B(_14355_), .Y(_14357_) );
	AOI21X1 AOI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_14357_), .B(_14348_), .C(_14344_), .Y(_14358_) );
	OAI21X1 OAI21X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_14358_), .B(_14353_), .C(_14342_), .Y(_14359_) );
	NAND3X1 NAND3X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_14359_), .B(_14352_), .C(_14341_), .Y(_14360_) );
	OAI21X1 OAI21X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_14358_), .B(_14353_), .C(_14343_), .Y(_14361_) );
	NAND3X1 NAND3X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_14342_), .B(_14351_), .C(_14350_), .Y(_14362_) );
	NAND3X1 NAND3X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_14340_), .B(_14361_), .C(_14362_), .Y(_14363_) );
	AOI21X1 AOI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_14089_), .B(_14086_), .C(_14091_), .Y(_14364_) );
	OAI21X1 OAI21X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_14364_), .B(_14079_), .C(_14092_), .Y(_14365_) );
	NAND3X1 NAND3X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_14365_), .B(_14363_), .C(_14360_), .Y(_14366_) );
	AOI21X1 AOI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_14362_), .B(_14361_), .C(_14340_), .Y(_14368_) );
	AOI21X1 AOI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_14352_), .B(_14359_), .C(_14341_), .Y(_14369_) );
	INVX1 INVX1_1926 ( .gnd(gnd), .vdd(vdd), .A(_14092_), .Y(_14370_) );
	AOI21X1 AOI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_14078_), .B(_14099_), .C(_14370_), .Y(_14371_) );
	OAI21X1 OAI21X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_14369_), .B(_14368_), .C(_14371_), .Y(_14372_) );
	NAND3X1 NAND3X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_14329_), .B(_14366_), .C(_14372_), .Y(_14373_) );
	NAND2X1 NAND2X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_14046_), .B(_14053_), .Y(_14374_) );
	NAND3X1 NAND3X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_14363_), .B(_14371_), .C(_14360_), .Y(_14375_) );
	OAI21X1 OAI21X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_14369_), .B(_14368_), .C(_14365_), .Y(_14376_) );
	NAND3X1 NAND3X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_14374_), .B(_14375_), .C(_14376_), .Y(_14377_) );
	NAND2X1 NAND2X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_14373_), .B(_14377_), .Y(_14379_) );
	AOI21X1 AOI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_14146_), .B(_14140_), .C(_14107_), .Y(_14380_) );
	OAI21X1 OAI21X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_14157_), .B(_14380_), .C(_14147_), .Y(_14381_) );
	NAND2X1 NAND2X1_2869 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf1), .B(aOperand_frameOut_16_bF_buf3), .Y(_14382_) );
	OAI21X1 OAI21X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_13773_), .B(_14382_), .C(_14086_), .Y(_14383_) );
	INVX1 INVX1_1927 ( .gnd(gnd), .vdd(vdd), .A(_14383_), .Y(_14384_) );
	NOR2X1 NOR2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf0), .B(_12233_), .Y(_14385_) );
	NAND2X1 NAND2X1_2870 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf0), .B(aOperand_frameOut_17_bF_buf0), .Y(_14386_) );
	INVX1 INVX1_1928 ( .gnd(gnd), .vdd(vdd), .A(_14386_), .Y(_14387_) );
	NAND2X1 NAND2X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_14083_), .B(_14387_), .Y(_14388_) );
	OAI21X1 OAI21X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf3), .B(_12708_), .C(_14382_), .Y(_14390_) );
	NAND3X1 NAND3X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_14385_), .B(_14390_), .C(_14388_), .Y(_14391_) );
	NAND2X1 NAND2X1_2872 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf1), .B(aOperand_frameOut_16_bF_buf2), .Y(_14392_) );
	OAI21X1 OAI21X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_14392_), .B(_14386_), .C(_14390_), .Y(_14393_) );
	OAI21X1 OAI21X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf3), .B(_12233_), .C(_14393_), .Y(_14394_) );
	AOI21X1 AOI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_14113_), .B(_14108_), .C(_14111_), .Y(_14395_) );
	INVX1 INVX1_1929 ( .gnd(gnd), .vdd(vdd), .A(_14395_), .Y(_14396_) );
	NAND3X1 NAND3X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_14391_), .B(_14394_), .C(_14396_), .Y(_14397_) );
	INVX1 INVX1_1930 ( .gnd(gnd), .vdd(vdd), .A(_14385_), .Y(_14398_) );
	NOR2X1 NOR2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_14398_), .B(_14393_), .Y(_14399_) );
	AOI21X1 AOI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_14388_), .B(_14390_), .C(_14385_), .Y(_14401_) );
	OAI21X1 OAI21X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_14401_), .B(_14399_), .C(_14395_), .Y(_14402_) );
	NAND3X1 NAND3X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_14384_), .B(_14397_), .C(_14402_), .Y(_14403_) );
	NAND3X1 NAND3X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_14395_), .B(_14391_), .C(_14394_), .Y(_14404_) );
	OAI21X1 OAI21X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_14401_), .B(_14399_), .C(_14396_), .Y(_14405_) );
	NAND3X1 NAND3X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_14383_), .B(_14404_), .C(_14405_), .Y(_14406_) );
	NAND2X1 NAND2X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_14403_), .B(_14406_), .Y(_14407_) );
	AOI21X1 AOI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_14129_), .B(_14133_), .C(_14119_), .Y(_14408_) );
	OAI21X1 OAI21X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_14408_), .B(_14143_), .C(_14134_), .Y(_14409_) );
	NOR2X1 NOR2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf2), .B(_13796_), .Y(_14410_) );
	INVX1 INVX1_1931 ( .gnd(gnd), .vdd(vdd), .A(_14410_), .Y(_14412_) );
	INVX1 INVX1_1932 ( .gnd(gnd), .vdd(vdd), .A(_14110_), .Y(_14413_) );
	NAND2X1 NAND2X1_2874 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .B(aOperand_frameOut_20_bF_buf2), .Y(_14414_) );
	INVX1 INVX1_1933 ( .gnd(gnd), .vdd(vdd), .A(_14414_), .Y(_14415_) );
	NAND2X1 NAND2X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_14413_), .B(_14415_), .Y(_14416_) );
	NAND2X1 NAND2X1_2876 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .B(aOperand_frameOut_20_bF_buf1), .Y(_14417_) );
	OAI21X1 OAI21X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_13224_), .C(_14417_), .Y(_14418_) );
	NAND3X1 NAND3X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_14418_), .B(_14416_), .C(_14412_), .Y(_14419_) );
	OAI21X1 OAI21X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_14110_), .B(_14414_), .C(_14418_), .Y(_14420_) );
	NAND2X1 NAND2X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_14410_), .B(_14420_), .Y(_14421_) );
	NAND2X1 NAND2X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_14419_), .B(_14421_), .Y(_14423_) );
	NOR2X1 NOR2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_14122_), .B(_14123_), .Y(_14424_) );
	OAI21X1 OAI21X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_14120_), .B(_14424_), .C(_14124_), .Y(_14425_) );
	NAND2X1 NAND2X1_2879 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf3), .B(aOperand_frameOut_21_bF_buf2), .Y(_14426_) );
	INVX1 INVX1_1934 ( .gnd(gnd), .vdd(vdd), .A(_14426_), .Y(_14427_) );
	AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(aOperand_frameOut_22_bF_buf0), .Y(_14428_) );
	AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_23_), .Y(_14429_) );
	NAND2X1 NAND2X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_14428_), .B(_14429_), .Y(_14430_) );
	NAND2X1 NAND2X1_2881 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(aOperand_frameOut_23_), .Y(_14431_) );
	OAI21X1 OAI21X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf1), .B(_14125_), .C(_14431_), .Y(_14432_) );
	NAND3X1 NAND3X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_14427_), .B(_14432_), .C(_14430_), .Y(_14434_) );
	OAI21X1 OAI21X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf0), .B(_14125_), .C(_14429_), .Y(_14435_) );
	INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_23_), .Y(_14436_) );
	OAI21X1 OAI21X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf4), .B(_14436_), .C(_14428_), .Y(_14437_) );
	NAND3X1 NAND3X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_14426_), .B(_14435_), .C(_14437_), .Y(_14438_) );
	NAND3X1 NAND3X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_14434_), .B(_14438_), .C(_14425_), .Y(_14439_) );
	AOI22X1 AOI22X1_340 ( .gnd(gnd), .vdd(vdd), .A(_13810_), .B(_14428_), .C(_14121_), .D(_14128_), .Y(_14440_) );
	AOI21X1 AOI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_14435_), .B(_14437_), .C(_14426_), .Y(_14441_) );
	AOI22X1 AOI22X1_341 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf2), .B(aOperand_frameOut_21_bF_buf1), .C(_14432_), .D(_14430_), .Y(_14442_) );
	OAI21X1 OAI21X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_14442_), .B(_14441_), .C(_14440_), .Y(_14443_) );
	NAND3X1 NAND3X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_14423_), .B(_14439_), .C(_14443_), .Y(_14445_) );
	AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_14421_), .B(_14419_), .Y(_14446_) );
	OAI21X1 OAI21X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_14442_), .B(_14441_), .C(_14425_), .Y(_14447_) );
	NAND3X1 NAND3X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_14440_), .B(_14434_), .C(_14438_), .Y(_14448_) );
	NAND3X1 NAND3X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_14448_), .B(_14447_), .C(_14446_), .Y(_14449_) );
	NAND3X1 NAND3X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_14445_), .B(_14409_), .C(_14449_), .Y(_14450_) );
	NOR3X1 NOR3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_14136_), .B(_14135_), .C(_14138_), .Y(_14451_) );
	AOI21X1 AOI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_14118_), .B(_14139_), .C(_14451_), .Y(_14452_) );
	AOI22X1 AOI22X1_342 ( .gnd(gnd), .vdd(vdd), .A(_14419_), .B(_14421_), .C(_14448_), .D(_14447_), .Y(_14453_) );
	AOI21X1 AOI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_14443_), .B(_14439_), .C(_14423_), .Y(_14454_) );
	OAI21X1 OAI21X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_14453_), .B(_14454_), .C(_14452_), .Y(_14456_) );
	NAND3X1 NAND3X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_14450_), .B(_14407_), .C(_14456_), .Y(_14457_) );
	AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_14403_), .B(_14406_), .Y(_14458_) );
	OAI21X1 OAI21X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_14453_), .B(_14454_), .C(_14409_), .Y(_14459_) );
	NAND3X1 NAND3X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_14445_), .B(_14452_), .C(_14449_), .Y(_14460_) );
	NAND3X1 NAND3X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_14460_), .B(_14459_), .C(_14458_), .Y(_14461_) );
	NAND3X1 NAND3X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_14381_), .B(_14457_), .C(_14461_), .Y(_14462_) );
	NOR3X1 NOR3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_14151_), .B(_14152_), .C(_14150_), .Y(_14463_) );
	AOI21X1 AOI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_14105_), .B(_14153_), .C(_14463_), .Y(_14464_) );
	AOI22X1 AOI22X1_343 ( .gnd(gnd), .vdd(vdd), .A(_14403_), .B(_14406_), .C(_14460_), .D(_14459_), .Y(_14465_) );
	AOI21X1 AOI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_14456_), .B(_14450_), .C(_14407_), .Y(_14467_) );
	OAI21X1 OAI21X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_14465_), .B(_14467_), .C(_14464_), .Y(_14468_) );
	NAND3X1 NAND3X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_14462_), .B(_14468_), .C(_14379_), .Y(_14469_) );
	NAND3X1 NAND3X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_14374_), .B(_14366_), .C(_14372_), .Y(_14470_) );
	NAND3X1 NAND3X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_14329_), .B(_14375_), .C(_14376_), .Y(_14471_) );
	NAND2X1 NAND2X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14471_), .Y(_14472_) );
	OAI21X1 OAI21X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_14465_), .B(_14467_), .C(_14381_), .Y(_14473_) );
	NAND3X1 NAND3X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_14457_), .B(_14461_), .C(_14464_), .Y(_14474_) );
	NAND3X1 NAND3X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_14473_), .B(_14474_), .C(_14472_), .Y(_14475_) );
	NAND3X1 NAND3X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_14469_), .B(_14475_), .C(_14328_), .Y(_14476_) );
	INVX1 INVX1_1935 ( .gnd(gnd), .vdd(vdd), .A(_14162_), .Y(_14478_) );
	AOI21X1 AOI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_14074_), .B(_14167_), .C(_14478_), .Y(_14479_) );
	AOI22X1 AOI22X1_344 ( .gnd(gnd), .vdd(vdd), .A(_14373_), .B(_14377_), .C(_14473_), .D(_14474_), .Y(_14480_) );
	AOI22X1 AOI22X1_345 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14471_), .C(_14462_), .D(_14468_), .Y(_14481_) );
	OAI21X1 OAI21X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_14481_), .B(_14480_), .C(_14479_), .Y(_14482_) );
	NAND3X1 NAND3X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_14476_), .B(_14482_), .C(_14326_), .Y(_14483_) );
	NAND3X1 NAND3X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_14321_), .B(_14314_), .C(_14319_), .Y(_14484_) );
	NAND3X1 NAND3X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_14248_), .B(_14324_), .C(_14322_), .Y(_14485_) );
	NAND2X1 NAND2X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_14484_), .B(_14485_), .Y(_14486_) );
	OAI21X1 OAI21X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_14481_), .B(_14480_), .C(_14328_), .Y(_14487_) );
	NAND3X1 NAND3X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_14469_), .B(_14475_), .C(_14479_), .Y(_14488_) );
	NAND3X1 NAND3X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_14487_), .B(_14488_), .C(_14486_), .Y(_14489_) );
	NAND3X1 NAND3X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_14483_), .B(_14489_), .C(_14247_), .Y(_14490_) );
	NOR3X1 NOR3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_14180_), .B(_14179_), .C(_14178_), .Y(_14491_) );
	AOI21X1 AOI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_14024_), .B(_14182_), .C(_14491_), .Y(_14492_) );
	AOI22X1 AOI22X1_346 ( .gnd(gnd), .vdd(vdd), .A(_14320_), .B(_14325_), .C(_14487_), .D(_14488_), .Y(_14493_) );
	AOI22X1 AOI22X1_347 ( .gnd(gnd), .vdd(vdd), .A(_14484_), .B(_14485_), .C(_14476_), .D(_14482_), .Y(_14494_) );
	OAI21X1 OAI21X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_14494_), .B(_14493_), .C(_14492_), .Y(_14495_) );
	NAND3X1 NAND3X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_14244_), .B(_14490_), .C(_14495_), .Y(_14496_) );
	INVX1 INVX1_1936 ( .gnd(gnd), .vdd(vdd), .A(_14240_), .Y(_14497_) );
	NAND2X1 NAND2X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_14497_), .B(_14241_), .Y(_14500_) );
	OR2X2 OR2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_14241_), .B(_14497_), .Y(_14501_) );
	NAND2X1 NAND2X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .B(_14501_), .Y(_14502_) );
	OAI21X1 OAI21X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_14494_), .B(_14493_), .C(_14247_), .Y(_14503_) );
	NAND3X1 NAND3X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_14483_), .B(_14489_), .C(_14492_), .Y(_14504_) );
	NAND3X1 NAND3X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_14502_), .B(_14503_), .C(_14504_), .Y(_14505_) );
	NAND3X1 NAND3X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14505_), .C(_14234_), .Y(_14506_) );
	NOR3X1 NOR3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_14195_), .B(_14194_), .C(_14193_), .Y(_14507_) );
	AOI21X1 AOI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_13937_), .B(_14196_), .C(_14507_), .Y(_14508_) );
	AOI22X1 AOI22X1_348 ( .gnd(gnd), .vdd(vdd), .A(_14242_), .B(_14243_), .C(_14503_), .D(_14504_), .Y(_14509_) );
	AOI22X1 AOI22X1_349 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .B(_14501_), .C(_14490_), .D(_14495_), .Y(_14511_) );
	OAI21X1 OAI21X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_14511_), .B(_14509_), .C(_14508_), .Y(_14512_) );
	NAND3X1 NAND3X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_14232_), .B(_14506_), .C(_14512_), .Y(_14513_) );
	OAI21X1 OAI21X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_14511_), .B(_14509_), .C(_14234_), .Y(_14514_) );
	NAND3X1 NAND3X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14505_), .C(_14508_), .Y(_14515_) );
	NAND3X1 NAND3X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_14198_), .B(_14514_), .C(_14515_), .Y(_14516_) );
	NAND3X1 NAND3X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_14513_), .B(_14516_), .C(_14231_), .Y(_14517_) );
	NOR3X1 NOR3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_14208_), .B(_14207_), .C(_14206_), .Y(_14518_) );
	AOI21X1 AOI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_13619_), .B(_14209_), .C(_14518_), .Y(_14519_) );
	AOI21X1 AOI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_14515_), .B(_14514_), .C(_14198_), .Y(_14520_) );
	AOI22X1 AOI22X1_350 ( .gnd(gnd), .vdd(vdd), .A(_13932_), .B(_13934_), .C(_14506_), .D(_14512_), .Y(_14522_) );
	OAI21X1 OAI21X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_14522_), .B(_14520_), .C(_14519_), .Y(_14523_) );
	NAND3X1 NAND3X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_14215_), .B(_14517_), .C(_14523_), .Y(_14524_) );
	AOI21X1 AOI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_14217_), .B(_14216_), .C(_13887_), .Y(_14525_) );
	OAI21X1 OAI21X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_14522_), .B(_14520_), .C(_14231_), .Y(_14526_) );
	NAND3X1 NAND3X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_14513_), .B(_14516_), .C(_14519_), .Y(_14527_) );
	NAND3X1 NAND3X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_14525_), .B(_14526_), .C(_14527_), .Y(_14528_) );
	NAND2X1 NAND2X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_14524_), .B(_14528_), .Y(_14529_) );
	XNOR2X1 XNOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_14229_), .B(_14529_), .Y(mulOut_23_) );
	AOI22X1 AOI22X1_351 ( .gnd(gnd), .vdd(vdd), .A(_14219_), .B(_14222_), .C(_14524_), .D(_14528_), .Y(_14530_) );
	NAND2X1 NAND2X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_13925_), .B(_14530_), .Y(_14531_) );
	NOR3X1 NOR3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_13321_), .B(_14531_), .C(_12331_), .Y(_14532_) );
	AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_13905_), .B(_13903_), .Y(_14533_) );
	NAND3X1 NAND3X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_14215_), .B(_14526_), .C(_14527_), .Y(_14534_) );
	NAND3X1 NAND3X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_14517_), .B(_14525_), .C(_14523_), .Y(_14535_) );
	NAND2X1 NAND2X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_14227_), .B(_14535_), .Y(_14536_) );
	AOI22X1 AOI22X1_352 ( .gnd(gnd), .vdd(vdd), .A(_14534_), .B(_14536_), .C(_14530_), .D(_14533_), .Y(_14537_) );
	OAI21X1 OAI21X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_14531_), .B(_13325_), .C(_14537_), .Y(_14538_) );
	NOR2X1 NOR2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_14538_), .B(_14532_), .Y(_14539_) );
	NAND2X1 NAND2X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_14506_), .B(_14513_), .Y(_14540_) );
	INVX1 INVX1_1937 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .Y(_14542_) );
	NAND2X1 NAND2X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_14490_), .B(_14496_), .Y(_14543_) );
	INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_24_), .Y(_14544_) );
	NOR2X1 NOR2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf3), .B(_14544_), .Y(_14545_) );
	NAND3X1 NAND3X1_3120 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf1), .B(adder_bOperand_23_), .C(_14251_), .Y(_14546_) );
	OAI21X1 OAI21X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_13944_), .B(_14250_), .C(_14546_), .Y(_14547_) );
	XOR2X1 XOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_14547_), .B(_14545_), .Y(_14548_) );
	OAI21X1 OAI21X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_14264_), .B(_14253_), .C(_14271_), .Y(_14549_) );
	NAND2X1 NAND2X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_14549_), .B(_14548_), .Y(_14550_) );
	OR2X2 OR2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_14548_), .B(_14549_), .Y(_14551_) );
	NAND2X1 NAND2X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_14550_), .B(_14551_), .Y(_14553_) );
	XOR2X1 XOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_14553_), .B(_14239_), .Y(_14554_) );
	NAND2X1 NAND2X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_14314_), .B(_14484_), .Y(_14555_) );
	NAND2X1 NAND2X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_14554_), .B(_14555_), .Y(_14556_) );
	OR2X2 OR2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_14555_), .B(_14554_), .Y(_14557_) );
	NAND2X1 NAND2X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .B(_14557_), .Y(_14558_) );
	INVX1 INVX1_1938 ( .gnd(gnd), .vdd(vdd), .A(_14558_), .Y(_14559_) );
	NAND2X1 NAND2X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_14476_), .B(_14483_), .Y(_14560_) );
	NAND2X1 NAND2X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_14300_), .B(_14306_), .Y(_14561_) );
	INVX1 INVX1_1939 ( .gnd(gnd), .vdd(vdd), .A(_14561_), .Y(_14562_) );
	INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_23_), .Y(_14564_) );
	NAND2X1 NAND2X1_2898 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(adder_bOperand_22_bF_buf1), .Y(_14565_) );
	INVX1 INVX1_1940 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_22_bF_buf0), .Y(_14566_) );
	NAND2X1 NAND2X1_2899 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf0), .B(adder_bOperand_21_bF_buf0), .Y(_14567_) );
	OAI21X1 OAI21X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf1), .B(_14566_), .C(_14567_), .Y(_14568_) );
	OAI21X1 OAI21X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_14250_), .B(_14565_), .C(_14568_), .Y(_14569_) );
	OAI21X1 OAI21X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_11874_), .B(_14564_), .C(_14569_), .Y(_14570_) );
	NAND2X1 NAND2X1_2900 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf0), .B(adder_bOperand_23_), .Y(_14571_) );
	OR2X2 OR2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_14569_), .B(_14571_), .Y(_14572_) );
	NAND2X1 NAND2X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_14570_), .B(_14572_), .Y(_14573_) );
	OAI21X1 OAI21X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_13949_), .B(_14258_), .C(_14262_), .Y(_14575_) );
	NAND2X1 NAND2X1_2902 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .B(adder_bOperand_20_bF_buf2), .Y(_14576_) );
	INVX1 INVX1_1941 ( .gnd(gnd), .vdd(vdd), .A(_14576_), .Y(_14577_) );
	NAND2X1 NAND2X1_2903 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf0), .B(adder_bOperand_19_bF_buf0), .Y(_14578_) );
	OAI21X1 OAI21X1_3120 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf2), .B(_13338_), .C(_14258_), .Y(_14579_) );
	OAI21X1 OAI21X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_14259_), .B(_14578_), .C(_14579_), .Y(_14580_) );
	XNOR2X1 XNOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .B(_14577_), .Y(_14581_) );
	NOR2X1 NOR2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_14581_), .B(_14575_), .Y(_14582_) );
	INVX1 INVX1_1942 ( .gnd(gnd), .vdd(vdd), .A(_13949_), .Y(_14583_) );
	INVX1 INVX1_1943 ( .gnd(gnd), .vdd(vdd), .A(_14258_), .Y(_14584_) );
	AOI21X1 AOI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_14583_), .B(_14584_), .C(_14265_), .Y(_14586_) );
	XNOR2X1 XNOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .B(_14576_), .Y(_14587_) );
	NOR2X1 NOR2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_14587_), .B(_14586_), .Y(_14588_) );
	OAI21X1 OAI21X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_14588_), .B(_14582_), .C(_14573_), .Y(_14589_) );
	INVX1 INVX1_1944 ( .gnd(gnd), .vdd(vdd), .A(_14573_), .Y(_14590_) );
	NAND2X1 NAND2X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_14587_), .B(_14586_), .Y(_14591_) );
	NAND2X1 NAND2X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_14581_), .B(_14575_), .Y(_14592_) );
	NAND3X1 NAND3X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_14590_), .B(_14591_), .C(_14592_), .Y(_14593_) );
	AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_14589_), .B(_14593_), .Y(_14594_) );
	NAND2X1 NAND2X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_14289_), .B(_14295_), .Y(_14595_) );
	OAI21X1 OAI21X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_14292_), .B(_14278_), .C(_14283_), .Y(_14597_) );
	NAND2X1 NAND2X1_2907 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf2), .B(adder_bOperand_17_bF_buf3), .Y(_14598_) );
	NAND2X1 NAND2X1_2908 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf1), .B(adder_bOperand_16_bF_buf2), .Y(_14599_) );
	OAI21X1 OAI21X1_3124 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf1), .B(_12131_), .C(_14277_), .Y(_14600_) );
	OAI21X1 OAI21X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_14282_), .B(_14599_), .C(_14600_), .Y(_14601_) );
	XOR2X1 XOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14598_), .Y(_14602_) );
	OAI21X1 OAI21X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_14336_), .B(_14337_), .C(_14335_), .Y(_14603_) );
	NAND2X1 NAND2X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_14603_), .B(_14602_), .Y(_14604_) );
	OAI21X1 OAI21X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_12566_), .C(_14601_), .Y(_14605_) );
	OR2X2 OR2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_14601_), .B(_14598_), .Y(_14606_) );
	NAND2X1 NAND2X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_14605_), .B(_14606_), .Y(_14608_) );
	AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_14335_), .B(_14332_), .Y(_14609_) );
	NAND2X1 NAND2X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_14609_), .B(_14608_), .Y(_14610_) );
	NAND3X1 NAND3X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_14597_), .B(_14604_), .C(_14610_), .Y(_14611_) );
	INVX1 INVX1_1945 ( .gnd(gnd), .vdd(vdd), .A(_14597_), .Y(_14612_) );
	NOR2X1 NOR2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_14609_), .B(_14608_), .Y(_14613_) );
	NOR2X1 NOR2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_14603_), .B(_14602_), .Y(_14614_) );
	OAI21X1 OAI21X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_14614_), .B(_14613_), .C(_14612_), .Y(_14615_) );
	NAND3X1 NAND3X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_14595_), .B(_14611_), .C(_14615_), .Y(_14616_) );
	AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_14295_), .B(_14289_), .Y(_14617_) );
	NAND2X1 NAND2X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_14602_), .B(_14609_), .Y(_14619_) );
	NAND2X1 NAND2X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_14603_), .B(_14608_), .Y(_14620_) );
	AOI21X1 AOI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_14620_), .B(_14619_), .C(_14612_), .Y(_14621_) );
	AOI21X1 AOI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_14610_), .B(_14604_), .C(_14597_), .Y(_14622_) );
	OAI21X1 OAI21X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_14621_), .B(_14622_), .C(_14617_), .Y(_14623_) );
	NAND3X1 NAND3X1_3124 ( .gnd(gnd), .vdd(vdd), .A(_14616_), .B(_14623_), .C(_14594_), .Y(_14624_) );
	NAND2X1 NAND2X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_14593_), .B(_14589_), .Y(_14625_) );
	OAI21X1 OAI21X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_14621_), .B(_14622_), .C(_14595_), .Y(_14626_) );
	NAND3X1 NAND3X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_14611_), .B(_14617_), .C(_14615_), .Y(_14627_) );
	NAND3X1 NAND3X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_14625_), .B(_14626_), .C(_14627_), .Y(_14628_) );
	NAND2X1 NAND2X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_14366_), .B(_14470_), .Y(_14630_) );
	NAND3X1 NAND3X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_14628_), .B(_14630_), .C(_14624_), .Y(_14631_) );
	AOI21X1 AOI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_14627_), .B(_14626_), .C(_14625_), .Y(_14632_) );
	AOI21X1 AOI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_14623_), .B(_14616_), .C(_14594_), .Y(_14633_) );
	AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14366_), .Y(_14634_) );
	OAI21X1 OAI21X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_14633_), .B(_14632_), .C(_14634_), .Y(_14635_) );
	NAND3X1 NAND3X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_14562_), .B(_14631_), .C(_14635_), .Y(_14636_) );
	NAND3X1 NAND3X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_14624_), .B(_14628_), .C(_14634_), .Y(_14637_) );
	OAI21X1 OAI21X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_14633_), .B(_14632_), .C(_14630_), .Y(_14638_) );
	NAND3X1 NAND3X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_14561_), .B(_14638_), .C(_14637_), .Y(_14639_) );
	NAND2X1 NAND2X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_14636_), .B(_14639_), .Y(_14641_) );
	NAND2X1 NAND2X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_14462_), .B(_14469_), .Y(_14642_) );
	NAND2X1 NAND2X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_14352_), .B(_14360_), .Y(_14643_) );
	INVX1 INVX1_1946 ( .gnd(gnd), .vdd(vdd), .A(_14643_), .Y(_14644_) );
	NOR2X1 NOR2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_12365_), .Y(_14645_) );
	NOR2X1 NOR2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf0), .B(_17319_), .Y(_14646_) );
	NAND2X1 NAND2X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .B(_14646_), .Y(_14647_) );
	OAI21X1 OAI21X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf3), .B(_17157_), .C(_14337_), .Y(_14648_) );
	NAND2X1 NAND2X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_14648_), .B(_14647_), .Y(_14649_) );
	XNOR2X1 XNOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_14649_), .B(_14645_), .Y(_14650_) );
	OAI21X1 OAI21X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_14346_), .B(_14349_), .C(_14357_), .Y(_14652_) );
	NOR2X1 NOR2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf3), .B(_11858_), .Y(_14653_) );
	NAND2X1 NAND2X1_2921 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf1), .B(aOperand_frameOut_15_bF_buf2), .Y(_14654_) );
	OAI21X1 OAI21X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf3), .B(_12233_), .C(_14347_), .Y(_14655_) );
	OAI21X1 OAI21X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_14354_), .B(_14654_), .C(_14655_), .Y(_14656_) );
	XNOR2X1 XNOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_14656_), .B(_14653_), .Y(_14657_) );
	NAND2X1 NAND2X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_14652_), .B(_14657_), .Y(_14658_) );
	INVX1 INVX1_1947 ( .gnd(gnd), .vdd(vdd), .A(_14652_), .Y(_14659_) );
	XOR2X1 XOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_14656_), .B(_14653_), .Y(_14660_) );
	NAND2X1 NAND2X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_14659_), .B(_14660_), .Y(_14661_) );
	NAND3X1 NAND3X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_14650_), .B(_14658_), .C(_14661_), .Y(_14663_) );
	INVX1 INVX1_1948 ( .gnd(gnd), .vdd(vdd), .A(_14645_), .Y(_14664_) );
	XNOR2X1 XNOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_14649_), .B(_14664_), .Y(_14665_) );
	NAND2X1 NAND2X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_14652_), .B(_14660_), .Y(_14666_) );
	NAND2X1 NAND2X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_14659_), .B(_14657_), .Y(_14667_) );
	NAND3X1 NAND3X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_14665_), .B(_14666_), .C(_14667_), .Y(_14668_) );
	NAND3X1 NAND3X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_14383_), .B(_14397_), .C(_14402_), .Y(_14669_) );
	NAND2X1 NAND2X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_14397_), .B(_14669_), .Y(_14670_) );
	NAND3X1 NAND3X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_14663_), .B(_14668_), .C(_14670_), .Y(_14671_) );
	AOI21X1 AOI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_14667_), .B(_14666_), .C(_14665_), .Y(_14672_) );
	AOI21X1 AOI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_14661_), .B(_14658_), .C(_14650_), .Y(_14674_) );
	AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_14669_), .B(_14397_), .Y(_14675_) );
	OAI21X1 OAI21X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_14672_), .B(_14674_), .C(_14675_), .Y(_14676_) );
	NAND3X1 NAND3X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_14644_), .B(_14671_), .C(_14676_), .Y(_14677_) );
	NAND3X1 NAND3X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_14663_), .B(_14668_), .C(_14675_), .Y(_14678_) );
	OAI21X1 OAI21X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_14672_), .B(_14674_), .C(_14670_), .Y(_14679_) );
	NAND3X1 NAND3X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_14643_), .B(_14679_), .C(_14678_), .Y(_14680_) );
	NAND2X1 NAND2X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_14677_), .B(_14680_), .Y(_14681_) );
	NAND2X1 NAND2X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_14450_), .B(_14457_), .Y(_14682_) );
	OAI21X1 OAI21X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_14398_), .B(_14393_), .C(_14388_), .Y(_14683_) );
	INVX1 INVX1_1949 ( .gnd(gnd), .vdd(vdd), .A(_14683_), .Y(_14685_) );
	NAND2X1 NAND2X1_2929 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf2), .B(aOperand_frameOut_16_bF_buf1), .Y(_14686_) );
	NAND2X1 NAND2X1_2930 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf0), .B(aOperand_frameOut_17_bF_buf4), .Y(_14687_) );
	NAND2X1 NAND2X1_2931 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(aOperand_frameOut_18_bF_buf3), .Y(_14688_) );
	NAND2X1 NAND2X1_2932 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(aOperand_frameOut_18_bF_buf2), .Y(_14689_) );
	OAI21X1 OAI21X1_3140 ( .gnd(gnd), .vdd(vdd), .A(_13830_), .B(_12708_), .C(_14689_), .Y(_14690_) );
	OAI21X1 OAI21X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_14687_), .B(_14688_), .C(_14690_), .Y(_14691_) );
	XOR2X1 XOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_14691_), .B(_14686_), .Y(_14692_) );
	OAI21X1 OAI21X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_14412_), .B(_14420_), .C(_14416_), .Y(_14693_) );
	NAND2X1 NAND2X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_14693_), .B(_14692_), .Y(_14694_) );
	NOR2X1 NOR2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_14686_), .B(_14691_), .Y(_14696_) );
	AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_14691_), .B(_14686_), .Y(_14697_) );
	INVX1 INVX1_1950 ( .gnd(gnd), .vdd(vdd), .A(_14693_), .Y(_14698_) );
	OAI21X1 OAI21X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_14696_), .B(_14697_), .C(_14698_), .Y(_14699_) );
	NAND3X1 NAND3X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_14685_), .B(_14694_), .C(_14699_), .Y(_14700_) );
	NAND2X1 NAND2X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_14698_), .B(_14692_), .Y(_14701_) );
	OAI21X1 OAI21X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_14696_), .B(_14697_), .C(_14693_), .Y(_14702_) );
	NAND3X1 NAND3X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_14683_), .B(_14702_), .C(_14701_), .Y(_14703_) );
	NAND2X1 NAND2X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_14703_), .B(_14700_), .Y(_14704_) );
	NAND2X1 NAND2X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_14434_), .B(_14438_), .Y(_14705_) );
	OAI21X1 OAI21X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_14440_), .B(_14705_), .C(_14445_), .Y(_14707_) );
	NOR2X1 NOR2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf1), .B(_13224_), .Y(_14708_) );
	NAND2X1 NAND2X1_2937 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf3), .B(aOperand_frameOut_21_bF_buf0), .Y(_14709_) );
	OAI21X1 OAI21X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf3), .B(_13812_), .C(_14414_), .Y(_14710_) );
	OAI21X1 OAI21X1_3147 ( .gnd(gnd), .vdd(vdd), .A(_14417_), .B(_14709_), .C(_14710_), .Y(_14711_) );
	XNOR2X1 XNOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_14711_), .B(_14708_), .Y(_14712_) );
	NAND2X1 NAND2X1_2938 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf4), .B(aOperand_frameOut_23_), .Y(_14713_) );
	INVX1 INVX1_1951 ( .gnd(gnd), .vdd(vdd), .A(_14713_), .Y(_14714_) );
	AOI22X1 AOI22X1_353 ( .gnd(gnd), .vdd(vdd), .A(_14714_), .B(_14123_), .C(_14427_), .D(_14432_), .Y(_14715_) );
	INVX1 INVX1_1952 ( .gnd(gnd), .vdd(vdd), .A(_14715_), .Y(_14716_) );
	NOR2X1 NOR2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_14125_), .Y(_14718_) );
	NAND2X1 NAND2X1_2939 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf3), .B(aOperand_frameOut_24_bF_buf2), .Y(_14719_) );
	INVX1 INVX1_1953 ( .gnd(gnd), .vdd(vdd), .A(_14719_), .Y(_14720_) );
	NAND2X1 NAND2X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_14429_), .B(_14720_), .Y(_14721_) );
	INVX1 INVX1_1954 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_24_bF_buf1), .Y(_14722_) );
	OAI21X1 OAI21X1_3148 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf3), .B(_14722_), .C(_14713_), .Y(_14723_) );
	NAND3X1 NAND3X1_3140 ( .gnd(gnd), .vdd(vdd), .A(_14718_), .B(_14723_), .C(_14721_), .Y(_14724_) );
	OAI21X1 OAI21X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_14431_), .B(_14719_), .C(_14723_), .Y(_14725_) );
	OAI21X1 OAI21X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_14125_), .C(_14725_), .Y(_14726_) );
	NAND3X1 NAND3X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_14724_), .B(_14726_), .C(_14716_), .Y(_14727_) );
	INVX1 INVX1_1955 ( .gnd(gnd), .vdd(vdd), .A(_14718_), .Y(_14729_) );
	NOR2X1 NOR2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_14729_), .B(_14725_), .Y(_14730_) );
	AOI21X1 AOI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_14721_), .B(_14723_), .C(_14718_), .Y(_14731_) );
	OAI21X1 OAI21X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_14731_), .B(_14730_), .C(_14715_), .Y(_14732_) );
	NAND3X1 NAND3X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_14712_), .B(_14727_), .C(_14732_), .Y(_14733_) );
	XOR2X1 XOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_14711_), .B(_14708_), .Y(_14734_) );
	OAI21X1 OAI21X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_14731_), .B(_14730_), .C(_14716_), .Y(_14735_) );
	NAND3X1 NAND3X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_14715_), .B(_14724_), .C(_14726_), .Y(_14736_) );
	NAND3X1 NAND3X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_14734_), .B(_14736_), .C(_14735_), .Y(_14737_) );
	NAND3X1 NAND3X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_14733_), .B(_14737_), .C(_14707_), .Y(_14738_) );
	NOR2X1 NOR2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_14440_), .B(_14705_), .Y(_14739_) );
	AOI21X1 AOI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_14423_), .B(_14443_), .C(_14739_), .Y(_14740_) );
	AOI21X1 AOI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_14735_), .B(_14736_), .C(_14734_), .Y(_14741_) );
	AOI21X1 AOI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_14732_), .B(_14727_), .C(_14712_), .Y(_14742_) );
	OAI21X1 OAI21X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_14741_), .B(_14742_), .C(_14740_), .Y(_14743_) );
	NAND3X1 NAND3X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_14704_), .B(_14743_), .C(_14738_), .Y(_14744_) );
	AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_14700_), .B(_14703_), .Y(_14745_) );
	NOR3X1 NOR3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_14740_), .B(_14741_), .C(_14742_), .Y(_14746_) );
	AOI21X1 AOI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_14733_), .B(_14737_), .C(_14707_), .Y(_14747_) );
	OAI21X1 OAI21X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_14747_), .B(_14746_), .C(_14745_), .Y(_14748_) );
	NAND3X1 NAND3X1_3147 ( .gnd(gnd), .vdd(vdd), .A(_14682_), .B(_14744_), .C(_14748_), .Y(_14750_) );
	AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_14457_), .B(_14450_), .Y(_14751_) );
	OAI21X1 OAI21X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_14741_), .B(_14742_), .C(_14707_), .Y(_14752_) );
	NAND3X1 NAND3X1_3148 ( .gnd(gnd), .vdd(vdd), .A(_14737_), .B(_14733_), .C(_14740_), .Y(_14753_) );
	AOI21X1 AOI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_14752_), .B(_14753_), .C(_14745_), .Y(_14754_) );
	AOI21X1 AOI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_14738_), .B(_14743_), .C(_14704_), .Y(_14755_) );
	OAI21X1 OAI21X1_3156 ( .gnd(gnd), .vdd(vdd), .A(_14755_), .B(_14754_), .C(_14751_), .Y(_14756_) );
	NAND3X1 NAND3X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_14750_), .B(_14756_), .C(_14681_), .Y(_14757_) );
	NAND3X1 NAND3X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_14643_), .B(_14671_), .C(_14676_), .Y(_14758_) );
	NAND3X1 NAND3X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_14644_), .B(_14679_), .C(_14678_), .Y(_14759_) );
	NAND2X1 NAND2X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_14758_), .B(_14759_), .Y(_14762_) );
	OAI21X1 OAI21X1_3157 ( .gnd(gnd), .vdd(vdd), .A(_14755_), .B(_14754_), .C(_14682_), .Y(_14763_) );
	NAND3X1 NAND3X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_14744_), .B(_14748_), .C(_14751_), .Y(_14764_) );
	NAND3X1 NAND3X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_14762_), .B(_14763_), .C(_14764_), .Y(_14765_) );
	NAND3X1 NAND3X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_14757_), .B(_14765_), .C(_14642_), .Y(_14766_) );
	AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_14469_), .B(_14462_), .Y(_14767_) );
	AOI21X1 AOI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_14764_), .B(_14763_), .C(_14762_), .Y(_14768_) );
	AOI21X1 AOI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_14756_), .B(_14750_), .C(_14681_), .Y(_14769_) );
	OAI21X1 OAI21X1_3158 ( .gnd(gnd), .vdd(vdd), .A(_14769_), .B(_14768_), .C(_14767_), .Y(_14770_) );
	NAND3X1 NAND3X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_14766_), .B(_14770_), .C(_14641_), .Y(_14771_) );
	NAND3X1 NAND3X1_3156 ( .gnd(gnd), .vdd(vdd), .A(_14561_), .B(_14631_), .C(_14635_), .Y(_14773_) );
	NAND3X1 NAND3X1_3157 ( .gnd(gnd), .vdd(vdd), .A(_14562_), .B(_14638_), .C(_14637_), .Y(_14774_) );
	NAND2X1 NAND2X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_14773_), .B(_14774_), .Y(_14775_) );
	OAI21X1 OAI21X1_3159 ( .gnd(gnd), .vdd(vdd), .A(_14769_), .B(_14768_), .C(_14642_), .Y(_14776_) );
	NAND3X1 NAND3X1_3158 ( .gnd(gnd), .vdd(vdd), .A(_14757_), .B(_14765_), .C(_14767_), .Y(_14777_) );
	NAND3X1 NAND3X1_3159 ( .gnd(gnd), .vdd(vdd), .A(_14776_), .B(_14777_), .C(_14775_), .Y(_14778_) );
	NAND3X1 NAND3X1_3160 ( .gnd(gnd), .vdd(vdd), .A(_14771_), .B(_14560_), .C(_14778_), .Y(_14779_) );
	AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_14483_), .B(_14476_), .Y(_14780_) );
	AOI21X1 AOI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_14777_), .B(_14776_), .C(_14775_), .Y(_14781_) );
	AOI21X1 AOI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_14770_), .B(_14766_), .C(_14641_), .Y(_14782_) );
	OAI21X1 OAI21X1_3160 ( .gnd(gnd), .vdd(vdd), .A(_14782_), .B(_14781_), .C(_14780_), .Y(_14784_) );
	NAND3X1 NAND3X1_3161 ( .gnd(gnd), .vdd(vdd), .A(_14559_), .B(_14779_), .C(_14784_), .Y(_14785_) );
	OAI21X1 OAI21X1_3161 ( .gnd(gnd), .vdd(vdd), .A(_14782_), .B(_14781_), .C(_14560_), .Y(_14786_) );
	NAND3X1 NAND3X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_14771_), .B(_14778_), .C(_14780_), .Y(_14787_) );
	NAND3X1 NAND3X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_14558_), .B(_14787_), .C(_14786_), .Y(_14788_) );
	NAND3X1 NAND3X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14785_), .C(_14788_), .Y(_14789_) );
	AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_14496_), .B(_14490_), .Y(_14790_) );
	AOI21X1 AOI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_14786_), .B(_14787_), .C(_14558_), .Y(_14791_) );
	AOI22X1 AOI22X1_354 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .B(_14557_), .C(_14779_), .D(_14784_), .Y(_14792_) );
	OAI21X1 OAI21X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_14792_), .B(_14791_), .C(_14790_), .Y(_14793_) );
	NAND3X1 NAND3X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_14542_), .B(_14789_), .C(_14793_), .Y(_14795_) );
	OAI21X1 OAI21X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_14792_), .B(_14791_), .C(_14543_), .Y(_14796_) );
	NAND3X1 NAND3X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_14785_), .B(_14788_), .C(_14790_), .Y(_14797_) );
	NAND3X1 NAND3X1_3167 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .B(_14797_), .C(_14796_), .Y(_14798_) );
	NAND3X1 NAND3X1_3168 ( .gnd(gnd), .vdd(vdd), .A(_14540_), .B(_14795_), .C(_14798_), .Y(_14799_) );
	AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_14513_), .B(_14506_), .Y(_14800_) );
	AOI21X1 AOI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_14796_), .B(_14797_), .C(_14500_), .Y(_14801_) );
	AOI22X1 AOI22X1_355 ( .gnd(gnd), .vdd(vdd), .A(_14497_), .B(_14241_), .C(_14789_), .D(_14793_), .Y(_14802_) );
	OAI21X1 OAI21X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_14802_), .B(_14801_), .C(_14800_), .Y(_14803_) );
	NAND3X1 NAND3X1_3169 ( .gnd(gnd), .vdd(vdd), .A(_14517_), .B(_14799_), .C(_14803_), .Y(_14804_) );
	INVX1 INVX1_1956 ( .gnd(gnd), .vdd(vdd), .A(_14517_), .Y(_14806_) );
	OAI21X1 OAI21X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_14802_), .B(_14801_), .C(_14540_), .Y(_14807_) );
	NAND3X1 NAND3X1_3170 ( .gnd(gnd), .vdd(vdd), .A(_14795_), .B(_14798_), .C(_14800_), .Y(_14808_) );
	NAND3X1 NAND3X1_3171 ( .gnd(gnd), .vdd(vdd), .A(_14806_), .B(_14808_), .C(_14807_), .Y(_14809_) );
	NAND2X1 NAND2X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_14804_), .B(_14809_), .Y(_14810_) );
	XNOR2X1 XNOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_14539_), .B(_14810_), .Y(mulOut_24_) );
	INVX1 INVX1_1957 ( .gnd(gnd), .vdd(vdd), .A(_14539_), .Y(_14811_) );
	AOI21X1 AOI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_14807_), .B(_14808_), .C(_14517_), .Y(_14812_) );
	AOI21X1 AOI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_14811_), .B(_14810_), .C(_14812_), .Y(_14813_) );
	AOI21X1 AOI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_14788_), .B(_14785_), .C(_14543_), .Y(_14814_) );
	OAI21X1 OAI21X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_14500_), .B(_14814_), .C(_14789_), .Y(_14816_) );
	INVX1 INVX1_1958 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .Y(_14817_) );
	AOI21X1 AOI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_14778_), .B(_14771_), .C(_14560_), .Y(_14818_) );
	OAI21X1 OAI21X1_3167 ( .gnd(gnd), .vdd(vdd), .A(_14558_), .B(_14818_), .C(_14779_), .Y(_14819_) );
	NAND2X1 NAND2X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_13945_), .B(_14236_), .Y(_14820_) );
	OR2X2 OR2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_14553_), .B(_14820_), .Y(_14821_) );
	NAND2X1 NAND2X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_14631_), .B(_14773_), .Y(_14822_) );
	NAND2X1 NAND2X1_2946 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf5), .B(adder_bOperand_25_), .Y(_14823_) );
	INVX1 INVX1_1959 ( .gnd(gnd), .vdd(vdd), .A(_14823_), .Y(_14824_) );
	NAND2X1 NAND2X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_14824_), .B(_14545_), .Y(_14825_) );
	INVX1 INVX1_1960 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_25_), .Y(_14827_) );
	NAND2X1 NAND2X1_2948 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf4), .B(adder_bOperand_24_), .Y(_14828_) );
	OAI21X1 OAI21X1_3168 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf2), .B(_14827_), .C(_14828_), .Y(_14829_) );
	AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .B(_14829_), .Y(_14830_) );
	OAI21X1 OAI21X1_3169 ( .gnd(gnd), .vdd(vdd), .A(_14250_), .B(_14565_), .C(_14572_), .Y(_14831_) );
	NOR2X1 NOR2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_14830_), .B(_14831_), .Y(_14832_) );
	NAND2X1 NAND2X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_14830_), .B(_14831_), .Y(_14833_) );
	INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(_14833_), .Y(_14834_) );
	NOR2X1 NOR2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_14832_), .B(_14834_), .Y(_14835_) );
	OAI21X1 OAI21X1_3170 ( .gnd(gnd), .vdd(vdd), .A(_14573_), .B(_14582_), .C(_14592_), .Y(_14836_) );
	NOR2X1 NOR2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_14836_), .B(_14835_), .Y(_14838_) );
	INVX1 INVX1_1961 ( .gnd(gnd), .vdd(vdd), .A(_14838_), .Y(_14839_) );
	NAND2X1 NAND2X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_14836_), .B(_14835_), .Y(_14840_) );
	NAND2X1 NAND2X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_14840_), .B(_14839_), .Y(_14841_) );
	NAND2X1 NAND2X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_14545_), .B(_14547_), .Y(_14842_) );
	NAND2X1 NAND2X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_14842_), .B(_14550_), .Y(_14843_) );
	XNOR2X1 XNOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_14841_), .B(_14843_), .Y(_14844_) );
	NAND2X1 NAND2X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_14844_), .B(_14822_), .Y(_14845_) );
	XOR2X1 XOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_14841_), .B(_14843_), .Y(_14846_) );
	NAND3X1 NAND3X1_3172 ( .gnd(gnd), .vdd(vdd), .A(_14631_), .B(_14773_), .C(_14846_), .Y(_14847_) );
	NAND3X1 NAND3X1_3173 ( .gnd(gnd), .vdd(vdd), .A(_14821_), .B(_14847_), .C(_14845_), .Y(_14849_) );
	INVX1 INVX1_1962 ( .gnd(gnd), .vdd(vdd), .A(_14821_), .Y(_14850_) );
	NAND3X1 NAND3X1_3174 ( .gnd(gnd), .vdd(vdd), .A(_14631_), .B(_14773_), .C(_14844_), .Y(_14851_) );
	NAND2X1 NAND2X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_14846_), .B(_14822_), .Y(_14852_) );
	NAND3X1 NAND3X1_3175 ( .gnd(gnd), .vdd(vdd), .A(_14850_), .B(_14851_), .C(_14852_), .Y(_14853_) );
	NAND2X1 NAND2X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_14849_), .B(_14853_), .Y(_14854_) );
	AOI21X1 AOI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_14765_), .B(_14757_), .C(_14642_), .Y(_14855_) );
	OAI21X1 OAI21X1_3171 ( .gnd(gnd), .vdd(vdd), .A(_14855_), .B(_14775_), .C(_14766_), .Y(_14856_) );
	NAND2X1 NAND2X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_14616_), .B(_14624_), .Y(_14857_) );
	NOR2X1 NOR2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf0), .B(_14564_), .Y(_14858_) );
	INVX1 INVX1_1963 ( .gnd(gnd), .vdd(vdd), .A(_14858_), .Y(_14860_) );
	NAND2X1 NAND2X1_2958 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf2), .B(adder_bOperand_22_bF_buf3), .Y(_14861_) );
	INVX1 INVX1_1964 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_21_bF_buf3), .Y(_14862_) );
	OAI21X1 OAI21X1_3172 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf3), .B(_14862_), .C(_14565_), .Y(_14863_) );
	OAI21X1 OAI21X1_3173 ( .gnd(gnd), .vdd(vdd), .A(_14567_), .B(_14861_), .C(_14863_), .Y(_14864_) );
	OR2X2 OR2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_14864_), .B(_14860_), .Y(_14865_) );
	OAI21X1 OAI21X1_3174 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf3), .B(_14564_), .C(_14864_), .Y(_14866_) );
	NAND2X1 NAND2X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_14866_), .B(_14865_), .Y(_14867_) );
	INVX1 INVX1_1965 ( .gnd(gnd), .vdd(vdd), .A(_14867_), .Y(_14868_) );
	OAI22X1 OAI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(_14259_), .B(_14578_), .C(_14576_), .D(_14580_), .Y(_14869_) );
	NOR2X1 NOR2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_13334_), .Y(_14871_) );
	NAND2X1 NAND2X1_2960 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf4), .B(adder_bOperand_18_bF_buf0), .Y(_14872_) );
	NAND2X1 NAND2X1_2961 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf1), .B(adder_bOperand_19_bF_buf3), .Y(_14873_) );
	NAND2X1 NAND2X1_2962 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf0), .B(adder_bOperand_18_bF_buf3), .Y(_14874_) );
	OAI21X1 OAI21X1_3175 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf1), .B(_13067_), .C(_14874_), .Y(_14875_) );
	OAI21X1 OAI21X1_3176 ( .gnd(gnd), .vdd(vdd), .A(_14872_), .B(_14873_), .C(_14875_), .Y(_14876_) );
	XNOR2X1 XNOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_14876_), .B(_14871_), .Y(_14877_) );
	NAND2X1 NAND2X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_14869_), .B(_14877_), .Y(_14878_) );
	INVX1 INVX1_1966 ( .gnd(gnd), .vdd(vdd), .A(_14869_), .Y(_14879_) );
	XOR2X1 XOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_14876_), .B(_14871_), .Y(_14880_) );
	NAND2X1 NAND2X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_14880_), .B(_14879_), .Y(_14882_) );
	NAND3X1 NAND3X1_3176 ( .gnd(gnd), .vdd(vdd), .A(_14878_), .B(_14882_), .C(_14868_), .Y(_14883_) );
	NAND2X1 NAND2X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_14869_), .B(_14880_), .Y(_14884_) );
	NAND2X1 NAND2X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_14877_), .B(_14879_), .Y(_14885_) );
	NAND3X1 NAND3X1_3177 ( .gnd(gnd), .vdd(vdd), .A(_14867_), .B(_14884_), .C(_14885_), .Y(_14886_) );
	AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_14883_), .B(_14886_), .Y(_14887_) );
	OAI21X1 OAI21X1_3177 ( .gnd(gnd), .vdd(vdd), .A(_14612_), .B(_14614_), .C(_14604_), .Y(_14888_) );
	NAND2X1 NAND2X1_2967 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf0), .B(adder_bOperand_15_bF_buf1), .Y(_14889_) );
	OR2X2 OR2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_14277_), .B(_14889_), .Y(_14890_) );
	OAI21X1 OAI21X1_3178 ( .gnd(gnd), .vdd(vdd), .A(_14598_), .B(_14601_), .C(_14890_), .Y(_14891_) );
	NAND2X1 NAND2X1_2968 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf0), .B(adder_bOperand_17_bF_buf2), .Y(_14893_) );
	NAND2X1 NAND2X1_2969 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf2), .B(adder_bOperand_16_bF_buf1), .Y(_14894_) );
	OAI21X1 OAI21X1_3179 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_12131_), .C(_14599_), .Y(_14895_) );
	OAI21X1 OAI21X1_3180 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14894_), .C(_14895_), .Y(_14896_) );
	XOR2X1 XOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .B(_14893_), .Y(_14897_) );
	AOI22X1 AOI22X1_356 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .B(_14646_), .C(_14645_), .D(_14648_), .Y(_14898_) );
	INVX1 INVX1_1967 ( .gnd(gnd), .vdd(vdd), .A(_14898_), .Y(_14899_) );
	NAND2X1 NAND2X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .B(_14897_), .Y(_14900_) );
	OAI21X1 OAI21X1_3181 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_12566_), .C(_14896_), .Y(_14901_) );
	OR2X2 OR2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_14896_), .B(_14893_), .Y(_14902_) );
	NAND2X1 NAND2X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_14901_), .B(_14902_), .Y(_14904_) );
	NAND2X1 NAND2X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_14898_), .B(_14904_), .Y(_14905_) );
	NAND3X1 NAND3X1_3178 ( .gnd(gnd), .vdd(vdd), .A(_14891_), .B(_14900_), .C(_14905_), .Y(_14906_) );
	INVX1 INVX1_1968 ( .gnd(gnd), .vdd(vdd), .A(_14891_), .Y(_14907_) );
	NAND2X1 NAND2X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_14898_), .B(_14897_), .Y(_14908_) );
	NAND2X1 NAND2X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .B(_14904_), .Y(_14909_) );
	NAND3X1 NAND3X1_3179 ( .gnd(gnd), .vdd(vdd), .A(_14907_), .B(_14908_), .C(_14909_), .Y(_14910_) );
	NAND3X1 NAND3X1_3180 ( .gnd(gnd), .vdd(vdd), .A(_14906_), .B(_14910_), .C(_14888_), .Y(_14911_) );
	AOI21X1 AOI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_14597_), .B(_14610_), .C(_14613_), .Y(_14912_) );
	AOI21X1 AOI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_14909_), .B(_14908_), .C(_14907_), .Y(_14913_) );
	AOI21X1 AOI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_14905_), .B(_14900_), .C(_14891_), .Y(_14915_) );
	OAI21X1 OAI21X1_3182 ( .gnd(gnd), .vdd(vdd), .A(_14915_), .B(_14913_), .C(_14912_), .Y(_14916_) );
	NAND3X1 NAND3X1_3181 ( .gnd(gnd), .vdd(vdd), .A(_14887_), .B(_14911_), .C(_14916_), .Y(_14917_) );
	NAND2X1 NAND2X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .B(_14883_), .Y(_14918_) );
	OAI21X1 OAI21X1_3183 ( .gnd(gnd), .vdd(vdd), .A(_14915_), .B(_14913_), .C(_14888_), .Y(_14919_) );
	NAND3X1 NAND3X1_3182 ( .gnd(gnd), .vdd(vdd), .A(_14906_), .B(_14910_), .C(_14912_), .Y(_14920_) );
	NAND3X1 NAND3X1_3183 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .B(_14920_), .C(_14919_), .Y(_14921_) );
	AOI21X1 AOI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_14663_), .B(_14668_), .C(_14670_), .Y(_14922_) );
	OAI21X1 OAI21X1_3184 ( .gnd(gnd), .vdd(vdd), .A(_14644_), .B(_14922_), .C(_14671_), .Y(_14923_) );
	AOI21X1 AOI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_14917_), .B(_14921_), .C(_14923_), .Y(_14924_) );
	NAND3X1 NAND3X1_3184 ( .gnd(gnd), .vdd(vdd), .A(_14923_), .B(_14917_), .C(_14921_), .Y(_14926_) );
	INVX1 INVX1_1969 ( .gnd(gnd), .vdd(vdd), .A(_14926_), .Y(_14927_) );
	OAI21X1 OAI21X1_3185 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .B(_14927_), .C(_14857_), .Y(_14928_) );
	AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_14624_), .B(_14616_), .Y(_14929_) );
	INVX1 INVX1_1970 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14930_) );
	NAND3X1 NAND3X1_3185 ( .gnd(gnd), .vdd(vdd), .A(_14926_), .B(_14929_), .C(_14930_), .Y(_14931_) );
	NAND2X1 NAND2X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_14931_), .B(_14928_), .Y(_14932_) );
	NAND2X1 NAND2X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_14750_), .B(_14757_), .Y(_14933_) );
	OAI21X1 OAI21X1_3186 ( .gnd(gnd), .vdd(vdd), .A(_14659_), .B(_14660_), .C(_14663_), .Y(_14934_) );
	NOR2X1 NOR2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_12365_), .Y(_14935_) );
	NAND2X1 NAND2X1_2978 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf1), .B(aOperand_frameOut_13_bF_buf2), .Y(_14937_) );
	INVX1 INVX1_1971 ( .gnd(gnd), .vdd(vdd), .A(_14937_), .Y(_14938_) );
	NAND2X1 NAND2X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14646_), .Y(_14939_) );
	OAI21X1 OAI21X1_3187 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf2), .B(_17319_), .C(_14937_), .Y(_14940_) );
	NAND2X1 NAND2X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_14939_), .Y(_14941_) );
	XNOR2X1 XNOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(_14935_), .Y(_14942_) );
	INVX1 INVX1_1972 ( .gnd(gnd), .vdd(vdd), .A(_14654_), .Y(_14943_) );
	AOI22X1 AOI22X1_357 ( .gnd(gnd), .vdd(vdd), .A(_14355_), .B(_14943_), .C(_14653_), .D(_14655_), .Y(_14944_) );
	INVX1 INVX1_1973 ( .gnd(gnd), .vdd(vdd), .A(_14944_), .Y(_14945_) );
	NAND2X1 NAND2X1_2981 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf3), .B(aOperand_frameOut_14_bF_buf4), .Y(_14946_) );
	NAND2X1 NAND2X1_2982 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf3), .B(aOperand_frameOut_15_bF_buf1), .Y(_14948_) );
	NAND2X1 NAND2X1_2983 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf0), .B(aOperand_frameOut_16_bF_buf0), .Y(_14949_) );
	NAND2X1 NAND2X1_2984 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf2), .B(aOperand_frameOut_16_bF_buf4), .Y(_14950_) );
	OAI21X1 OAI21X1_3188 ( .gnd(gnd), .vdd(vdd), .A(_16887_), .B(_12233_), .C(_14950_), .Y(_14951_) );
	OAI21X1 OAI21X1_3189 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14949_), .C(_14951_), .Y(_14952_) );
	XOR2X1 XOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .B(_14946_), .Y(_14953_) );
	NAND2X1 NAND2X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .B(_14953_), .Y(_14954_) );
	NOR2X1 NOR2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_14946_), .B(_14952_), .Y(_14955_) );
	AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .B(_14946_), .Y(_14956_) );
	OAI21X1 OAI21X1_3190 ( .gnd(gnd), .vdd(vdd), .A(_14955_), .B(_14956_), .C(_14944_), .Y(_14957_) );
	NAND3X1 NAND3X1_3186 ( .gnd(gnd), .vdd(vdd), .A(_14957_), .B(_14942_), .C(_14954_), .Y(_14959_) );
	INVX1 INVX1_1974 ( .gnd(gnd), .vdd(vdd), .A(_14935_), .Y(_14960_) );
	XNOR2X1 XNOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(_14960_), .Y(_14961_) );
	OAI21X1 OAI21X1_3191 ( .gnd(gnd), .vdd(vdd), .A(_14955_), .B(_14956_), .C(_14945_), .Y(_14962_) );
	NAND2X1 NAND2X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_14944_), .B(_14953_), .Y(_14963_) );
	NAND3X1 NAND3X1_3187 ( .gnd(gnd), .vdd(vdd), .A(_14961_), .B(_14962_), .C(_14963_), .Y(_14964_) );
	NOR2X1 NOR2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_14693_), .B(_14692_), .Y(_14965_) );
	OAI21X1 OAI21X1_3192 ( .gnd(gnd), .vdd(vdd), .A(_14685_), .B(_14965_), .C(_14694_), .Y(_14966_) );
	NAND3X1 NAND3X1_3188 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14964_), .C(_14966_), .Y(_14967_) );
	AOI21X1 AOI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_14963_), .B(_14962_), .C(_14961_), .Y(_14968_) );
	AOI21X1 AOI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14957_), .C(_14942_), .Y(_14970_) );
	AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_14692_), .B(_14693_), .Y(_14971_) );
	AOI21X1 AOI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_14683_), .B(_14699_), .C(_14971_), .Y(_14972_) );
	OAI21X1 OAI21X1_3193 ( .gnd(gnd), .vdd(vdd), .A(_14970_), .B(_14968_), .C(_14972_), .Y(_14973_) );
	NAND3X1 NAND3X1_3189 ( .gnd(gnd), .vdd(vdd), .A(_14934_), .B(_14967_), .C(_14973_), .Y(_14974_) );
	INVX1 INVX1_1975 ( .gnd(gnd), .vdd(vdd), .A(_14934_), .Y(_14975_) );
	NAND3X1 NAND3X1_3190 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14964_), .C(_14972_), .Y(_14976_) );
	OAI21X1 OAI21X1_3194 ( .gnd(gnd), .vdd(vdd), .A(_14968_), .B(_14970_), .C(_14966_), .Y(_14977_) );
	NAND3X1 NAND3X1_3191 ( .gnd(gnd), .vdd(vdd), .A(_14976_), .B(_14977_), .C(_14975_), .Y(_14978_) );
	AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_14978_), .B(_14974_), .Y(_14979_) );
	AOI21X1 AOI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_14704_), .B(_14743_), .C(_14746_), .Y(_14981_) );
	OAI22X1 OAI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(_14687_), .B(_14688_), .C(_14686_), .D(_14691_), .Y(_14982_) );
	OAI21X1 OAI21X1_3195 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf2), .B(_13224_), .C(_14688_), .Y(_14983_) );
	NAND2X1 NAND2X1_2987 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf4), .B(aOperand_frameOut_19_bF_buf4), .Y(_14984_) );
	OAI21X1 OAI21X1_3196 ( .gnd(gnd), .vdd(vdd), .A(_14689_), .B(_14984_), .C(_14983_), .Y(_14985_) );
	OAI21X1 OAI21X1_3197 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf2), .B(_12708_), .C(_14985_), .Y(_14986_) );
	NOR2X1 NOR2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf1), .B(_12708_), .Y(_14987_) );
	NOR2X1 NOR2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_14689_), .B(_14984_), .Y(_14988_) );
	INVX1 INVX1_1976 ( .gnd(gnd), .vdd(vdd), .A(_14988_), .Y(_14989_) );
	NAND3X1 NAND3X1_3192 ( .gnd(gnd), .vdd(vdd), .A(_14987_), .B(_14983_), .C(_14989_), .Y(_14990_) );
	NAND2X1 NAND2X1_2988 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf3), .B(aOperand_frameOut_21_bF_buf4), .Y(_14992_) );
	NOR2X1 NOR2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_14414_), .B(_14992_), .Y(_14993_) );
	AOI21X1 AOI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_14710_), .B(_14708_), .C(_14993_), .Y(_14994_) );
	INVX1 INVX1_1977 ( .gnd(gnd), .vdd(vdd), .A(_14994_), .Y(_14995_) );
	NAND3X1 NAND3X1_3193 ( .gnd(gnd), .vdd(vdd), .A(_14990_), .B(_14986_), .C(_14995_), .Y(_14996_) );
	AOI21X1 AOI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_14989_), .B(_14983_), .C(_14987_), .Y(_14997_) );
	INVX1 INVX1_1978 ( .gnd(gnd), .vdd(vdd), .A(_14987_), .Y(_14998_) );
	NOR2X1 NOR2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_14998_), .B(_14985_), .Y(_14999_) );
	OAI21X1 OAI21X1_3198 ( .gnd(gnd), .vdd(vdd), .A(_14999_), .B(_14997_), .C(_14994_), .Y(_15000_) );
	NAND3X1 NAND3X1_3194 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14996_), .C(_15000_), .Y(_15001_) );
	INVX1 INVX1_1979 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .Y(_15003_) );
	NAND3X1 NAND3X1_3195 ( .gnd(gnd), .vdd(vdd), .A(_14994_), .B(_14990_), .C(_14986_), .Y(_15004_) );
	OAI21X1 OAI21X1_3199 ( .gnd(gnd), .vdd(vdd), .A(_14999_), .B(_14997_), .C(_14995_), .Y(_15005_) );
	NAND3X1 NAND3X1_3196 ( .gnd(gnd), .vdd(vdd), .A(_15004_), .B(_15003_), .C(_15005_), .Y(_15006_) );
	AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_15001_), .B(_15006_), .Y(_15007_) );
	INVX1 INVX1_1980 ( .gnd(gnd), .vdd(vdd), .A(_14727_), .Y(_15008_) );
	AOI21X1 AOI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_14712_), .B(_14732_), .C(_15008_), .Y(_15009_) );
	NOR2X1 NOR2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf0), .B(_13514_), .Y(_15010_) );
	INVX1 INVX1_1981 ( .gnd(gnd), .vdd(vdd), .A(_15010_), .Y(_15011_) );
	NAND2X1 NAND2X1_2989 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf2), .B(aOperand_frameOut_22_bF_buf3), .Y(_15012_) );
	NAND2X1 NAND2X1_2990 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf2), .B(aOperand_frameOut_22_bF_buf2), .Y(_15014_) );
	OAI21X1 OAI21X1_3200 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_13812_), .C(_15014_), .Y(_15015_) );
	OAI21X1 OAI21X1_3201 ( .gnd(gnd), .vdd(vdd), .A(_14992_), .B(_15012_), .C(_15015_), .Y(_15016_) );
	OR2X2 OR2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_15016_), .B(_15011_), .Y(_15017_) );
	OAI21X1 OAI21X1_3202 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf3), .B(_13514_), .C(_15016_), .Y(_15018_) );
	NAND2X1 NAND2X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .B(_15017_), .Y(_15019_) );
	AOI22X1 AOI22X1_358 ( .gnd(gnd), .vdd(vdd), .A(_14720_), .B(_14429_), .C(_14718_), .D(_14723_), .Y(_15020_) );
	INVX1 INVX1_1982 ( .gnd(gnd), .vdd(vdd), .A(_15020_), .Y(_15021_) );
	NOR2X1 NOR2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_14436_), .Y(_15022_) );
	INVX1 INVX1_1983 ( .gnd(gnd), .vdd(vdd), .A(_15022_), .Y(_15023_) );
	NAND2X1 NAND2X1_2992 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf0), .B(aOperand_frameOut_24_bF_buf0), .Y(_15025_) );
	NAND2X1 NAND2X1_2993 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf2), .B(aOperand_frameOut_25_bF_buf3), .Y(_15026_) );
	INVX1 INVX1_1984 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_25_bF_buf2), .Y(_15027_) );
	OAI21X1 OAI21X1_3203 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf2), .B(_15027_), .C(_14719_), .Y(_15028_) );
	OAI21X1 OAI21X1_3204 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .B(_15026_), .C(_15028_), .Y(_15029_) );
	NOR2X1 NOR2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_15023_), .B(_15029_), .Y(_15030_) );
	INVX1 INVX1_1985 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .Y(_15031_) );
	INVX1 INVX1_1986 ( .gnd(gnd), .vdd(vdd), .A(_15026_), .Y(_15032_) );
	NAND2X1 NAND2X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_15031_), .B(_15032_), .Y(_15033_) );
	AOI21X1 AOI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_15028_), .C(_15022_), .Y(_15034_) );
	OAI21X1 OAI21X1_3205 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_15030_), .C(_15021_), .Y(_15036_) );
	NAND3X1 NAND3X1_3197 ( .gnd(gnd), .vdd(vdd), .A(_15022_), .B(_15028_), .C(_15033_), .Y(_15037_) );
	OAI21X1 OAI21X1_3206 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_14436_), .C(_15029_), .Y(_15038_) );
	NAND3X1 NAND3X1_3198 ( .gnd(gnd), .vdd(vdd), .A(_15020_), .B(_15037_), .C(_15038_), .Y(_15039_) );
	AOI21X1 AOI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_15036_), .B(_15039_), .C(_15019_), .Y(_15040_) );
	XNOR2X1 XNOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_15016_), .B(_15010_), .Y(_15041_) );
	NAND3X1 NAND3X1_3199 ( .gnd(gnd), .vdd(vdd), .A(_15037_), .B(_15038_), .C(_15021_), .Y(_15042_) );
	OAI21X1 OAI21X1_3207 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_15030_), .C(_15020_), .Y(_15043_) );
	AOI21X1 AOI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_15043_), .B(_15042_), .C(_15041_), .Y(_15044_) );
	OAI21X1 OAI21X1_3208 ( .gnd(gnd), .vdd(vdd), .A(_15040_), .B(_15044_), .C(_15009_), .Y(_15045_) );
	AOI21X1 AOI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_14726_), .B(_14724_), .C(_14716_), .Y(_15047_) );
	OAI21X1 OAI21X1_3209 ( .gnd(gnd), .vdd(vdd), .A(_14734_), .B(_15047_), .C(_14727_), .Y(_15048_) );
	NAND3X1 NAND3X1_3200 ( .gnd(gnd), .vdd(vdd), .A(_15041_), .B(_15042_), .C(_15043_), .Y(_15049_) );
	NAND3X1 NAND3X1_3201 ( .gnd(gnd), .vdd(vdd), .A(_15039_), .B(_15019_), .C(_15036_), .Y(_15050_) );
	NAND3X1 NAND3X1_3202 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .B(_15050_), .C(_15048_), .Y(_15051_) );
	AOI21X1 AOI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_15045_), .B(_15051_), .C(_15007_), .Y(_15052_) );
	NAND3X1 NAND3X1_3203 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .B(_15051_), .C(_15045_), .Y(_15053_) );
	INVX1 INVX1_1987 ( .gnd(gnd), .vdd(vdd), .A(_15053_), .Y(_15054_) );
	OAI21X1 OAI21X1_3210 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .B(_15054_), .C(_14981_), .Y(_15055_) );
	OAI21X1 OAI21X1_3211 ( .gnd(gnd), .vdd(vdd), .A(_14747_), .B(_14745_), .C(_14738_), .Y(_15056_) );
	INVX1 INVX1_1988 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .Y(_15058_) );
	AOI21X1 AOI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_15050_), .B(_15049_), .C(_15048_), .Y(_15059_) );
	INVX1 INVX1_1989 ( .gnd(gnd), .vdd(vdd), .A(_15051_), .Y(_15060_) );
	OAI21X1 OAI21X1_3212 ( .gnd(gnd), .vdd(vdd), .A(_15059_), .B(_15060_), .C(_15058_), .Y(_15061_) );
	NAND3X1 NAND3X1_3204 ( .gnd(gnd), .vdd(vdd), .A(_15053_), .B(_15056_), .C(_15061_), .Y(_15062_) );
	NAND3X1 NAND3X1_3205 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .B(_15055_), .C(_14979_), .Y(_15063_) );
	NAND2X1 NAND2X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14978_), .Y(_15064_) );
	AOI21X1 AOI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_15061_), .B(_15053_), .C(_15056_), .Y(_15065_) );
	NOR3X1 NOR3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_15052_), .C(_15054_), .Y(_15066_) );
	OAI21X1 OAI21X1_3213 ( .gnd(gnd), .vdd(vdd), .A(_15065_), .B(_15066_), .C(_15064_), .Y(_15067_) );
	NAND3X1 NAND3X1_3206 ( .gnd(gnd), .vdd(vdd), .A(_15063_), .B(_15067_), .C(_14933_), .Y(_15069_) );
	NOR3X1 NOR3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_14755_), .B(_14754_), .C(_14751_), .Y(_15070_) );
	AOI21X1 AOI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_14681_), .B(_14756_), .C(_15070_), .Y(_15071_) );
	NOR3X1 NOR3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_15064_), .B(_15065_), .C(_15066_), .Y(_15072_) );
	AOI21X1 AOI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .B(_15062_), .C(_14979_), .Y(_15073_) );
	OAI21X1 OAI21X1_3214 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_15072_), .C(_15071_), .Y(_15074_) );
	NAND3X1 NAND3X1_3207 ( .gnd(gnd), .vdd(vdd), .A(_15069_), .B(_14932_), .C(_15074_), .Y(_15075_) );
	NAND3X1 NAND3X1_3208 ( .gnd(gnd), .vdd(vdd), .A(_14857_), .B(_14926_), .C(_14930_), .Y(_15076_) );
	OAI21X1 OAI21X1_3215 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .B(_14927_), .C(_14929_), .Y(_15077_) );
	NAND2X1 NAND2X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_15076_), .B(_15077_), .Y(_15078_) );
	OAI21X1 OAI21X1_3216 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_15072_), .C(_14933_), .Y(_15080_) );
	NAND3X1 NAND3X1_3209 ( .gnd(gnd), .vdd(vdd), .A(_15071_), .B(_15063_), .C(_15067_), .Y(_15081_) );
	NAND3X1 NAND3X1_3210 ( .gnd(gnd), .vdd(vdd), .A(_15081_), .B(_15078_), .C(_15080_), .Y(_15082_) );
	NAND3X1 NAND3X1_3211 ( .gnd(gnd), .vdd(vdd), .A(_14856_), .B(_15082_), .C(_15075_), .Y(_15083_) );
	INVX1 INVX1_1990 ( .gnd(gnd), .vdd(vdd), .A(_14766_), .Y(_15084_) );
	AOI21X1 AOI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_14641_), .B(_14770_), .C(_15084_), .Y(_15085_) );
	AOI22X1 AOI22X1_359 ( .gnd(gnd), .vdd(vdd), .A(_14928_), .B(_14931_), .C(_15081_), .D(_15080_), .Y(_15086_) );
	AOI21X1 AOI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .B(_15069_), .C(_14932_), .Y(_15087_) );
	OAI21X1 OAI21X1_3217 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .B(_15087_), .C(_15085_), .Y(_15088_) );
	NAND3X1 NAND3X1_3212 ( .gnd(gnd), .vdd(vdd), .A(_14854_), .B(_15083_), .C(_15088_), .Y(_15089_) );
	NAND3X1 NAND3X1_3213 ( .gnd(gnd), .vdd(vdd), .A(_14821_), .B(_14851_), .C(_14852_), .Y(_15091_) );
	NAND3X1 NAND3X1_3214 ( .gnd(gnd), .vdd(vdd), .A(_14850_), .B(_14847_), .C(_14845_), .Y(_15092_) );
	NAND2X1 NAND2X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_15091_), .B(_15092_), .Y(_15093_) );
	OAI21X1 OAI21X1_3218 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .B(_15087_), .C(_14856_), .Y(_15094_) );
	NAND3X1 NAND3X1_3215 ( .gnd(gnd), .vdd(vdd), .A(_15085_), .B(_15082_), .C(_15075_), .Y(_15095_) );
	NAND3X1 NAND3X1_3216 ( .gnd(gnd), .vdd(vdd), .A(_15093_), .B(_15095_), .C(_15094_), .Y(_15096_) );
	NAND3X1 NAND3X1_3217 ( .gnd(gnd), .vdd(vdd), .A(_14819_), .B(_15096_), .C(_15089_), .Y(_15097_) );
	INVX1 INVX1_1991 ( .gnd(gnd), .vdd(vdd), .A(_14779_), .Y(_15098_) );
	AOI21X1 AOI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_14559_), .B(_14784_), .C(_15098_), .Y(_15099_) );
	AOI21X1 AOI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_15094_), .B(_15095_), .C(_15093_), .Y(_15100_) );
	AOI21X1 AOI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_15088_), .B(_15083_), .C(_14854_), .Y(_15102_) );
	OAI21X1 OAI21X1_3219 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .B(_15102_), .C(_15099_), .Y(_15103_) );
	NAND3X1 NAND3X1_3218 ( .gnd(gnd), .vdd(vdd), .A(_14817_), .B(_15097_), .C(_15103_), .Y(_15104_) );
	OAI21X1 OAI21X1_3220 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .B(_15102_), .C(_14819_), .Y(_15105_) );
	NAND3X1 NAND3X1_3219 ( .gnd(gnd), .vdd(vdd), .A(_15089_), .B(_15096_), .C(_15099_), .Y(_15106_) );
	NAND3X1 NAND3X1_3220 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .B(_15106_), .C(_15105_), .Y(_15107_) );
	NAND3X1 NAND3X1_3221 ( .gnd(gnd), .vdd(vdd), .A(_14816_), .B(_15104_), .C(_15107_), .Y(_15108_) );
	INVX1 INVX1_1992 ( .gnd(gnd), .vdd(vdd), .A(_14789_), .Y(_15109_) );
	AOI21X1 AOI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_14542_), .B(_14793_), .C(_15109_), .Y(_15110_) );
	AOI21X1 AOI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_15105_), .B(_15106_), .C(_14556_), .Y(_15111_) );
	AOI22X1 AOI22X1_360 ( .gnd(gnd), .vdd(vdd), .A(_14554_), .B(_14555_), .C(_15097_), .D(_15103_), .Y(_15113_) );
	OAI21X1 OAI21X1_3221 ( .gnd(gnd), .vdd(vdd), .A(_15113_), .B(_15111_), .C(_15110_), .Y(_15114_) );
	NAND3X1 NAND3X1_3222 ( .gnd(gnd), .vdd(vdd), .A(_14799_), .B(_15108_), .C(_15114_), .Y(_15115_) );
	INVX1 INVX1_1993 ( .gnd(gnd), .vdd(vdd), .A(_14799_), .Y(_15116_) );
	OAI21X1 OAI21X1_3222 ( .gnd(gnd), .vdd(vdd), .A(_15113_), .B(_15111_), .C(_14816_), .Y(_15117_) );
	NAND3X1 NAND3X1_3223 ( .gnd(gnd), .vdd(vdd), .A(_15110_), .B(_15104_), .C(_15107_), .Y(_15118_) );
	NAND3X1 NAND3X1_3224 ( .gnd(gnd), .vdd(vdd), .A(_15118_), .B(_15116_), .C(_15117_), .Y(_15119_) );
	NAND2X1 NAND2X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_15115_), .B(_15119_), .Y(_15120_) );
	XNOR2X1 XNOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_14813_), .B(_15120_), .Y(mulOut_25_) );
	NAND3X1 NAND3X1_3225 ( .gnd(gnd), .vdd(vdd), .A(_15108_), .B(_15116_), .C(_15114_), .Y(_15121_) );
	NAND3X1 NAND3X1_3226 ( .gnd(gnd), .vdd(vdd), .A(_14799_), .B(_15118_), .C(_15117_), .Y(_15123_) );
	NAND2X1 NAND2X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_14812_), .B(_15123_), .Y(_15124_) );
	AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_15124_), .B(_15121_), .Y(_15125_) );
	NAND3X1 NAND3X1_3227 ( .gnd(gnd), .vdd(vdd), .A(_15121_), .B(_15123_), .C(_14810_), .Y(_15126_) );
	OAI21X1 OAI21X1_3223 ( .gnd(gnd), .vdd(vdd), .A(_15126_), .B(_14539_), .C(_15125_), .Y(_15127_) );
	AOI21X1 AOI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_15089_), .B(_15096_), .C(_14819_), .Y(_15128_) );
	OAI21X1 OAI21X1_3224 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .B(_15128_), .C(_15097_), .Y(_15129_) );
	NAND2X1 NAND2X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_14845_), .B(_15092_), .Y(_15130_) );
	AOI21X1 AOI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_15075_), .B(_15082_), .C(_14856_), .Y(_15131_) );
	OAI21X1 OAI21X1_3225 ( .gnd(gnd), .vdd(vdd), .A(_15093_), .B(_15131_), .C(_15083_), .Y(_15132_) );
	NOR2X1 NOR2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_14550_), .B(_14841_), .Y(_15134_) );
	INVX1 INVX1_1994 ( .gnd(gnd), .vdd(vdd), .A(_14825_), .Y(_15135_) );
	NAND2X1 NAND2X1_3001 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf0), .B(adder_bOperand_26_), .Y(_15136_) );
	NAND2X1 NAND2X1_3002 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf3), .B(adder_bOperand_25_), .Y(_15137_) );
	OAI21X1 OAI21X1_3226 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf2), .B(_14544_), .C(_14823_), .Y(_15138_) );
	OAI21X1 OAI21X1_3227 ( .gnd(gnd), .vdd(vdd), .A(_14828_), .B(_15137_), .C(_15138_), .Y(_15139_) );
	XOR2X1 XOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_15139_), .B(_15136_), .Y(_15140_) );
	NAND2X1 NAND2X1_3003 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf1), .B(adder_bOperand_21_bF_buf2), .Y(_15141_) );
	NOR2X1 NOR2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_14565_), .B(_15141_), .Y(_15142_) );
	AOI21X1 AOI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_14863_), .B(_14858_), .C(_15142_), .Y(_15143_) );
	INVX1 INVX1_1995 ( .gnd(gnd), .vdd(vdd), .A(_15143_), .Y(_15145_) );
	NAND2X1 NAND2X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_15145_), .B(_15140_), .Y(_15146_) );
	XNOR2X1 XNOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_15139_), .B(_15136_), .Y(_15147_) );
	NAND2X1 NAND2X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_15143_), .B(_15147_), .Y(_15148_) );
	AOI21X1 AOI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_15146_), .B(_15148_), .C(_15135_), .Y(_15149_) );
	INVX1 INVX1_1996 ( .gnd(gnd), .vdd(vdd), .A(_15149_), .Y(_15150_) );
	NAND3X1 NAND3X1_3228 ( .gnd(gnd), .vdd(vdd), .A(_15135_), .B(_15148_), .C(_15146_), .Y(_15151_) );
	INVX1 INVX1_1997 ( .gnd(gnd), .vdd(vdd), .A(_14878_), .Y(_15152_) );
	AOI21X1 AOI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_14868_), .B(_14882_), .C(_15152_), .Y(_15153_) );
	NAND3X1 NAND3X1_3229 ( .gnd(gnd), .vdd(vdd), .A(_15151_), .B(_15153_), .C(_15150_), .Y(_15154_) );
	INVX1 INVX1_1998 ( .gnd(gnd), .vdd(vdd), .A(_15151_), .Y(_15156_) );
	OAI21X1 OAI21X1_3228 ( .gnd(gnd), .vdd(vdd), .A(_14879_), .B(_14880_), .C(_14883_), .Y(_15157_) );
	OAI21X1 OAI21X1_3229 ( .gnd(gnd), .vdd(vdd), .A(_15149_), .B(_15156_), .C(_15157_), .Y(_15158_) );
	AOI21X1 AOI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_15158_), .B(_15154_), .C(_14833_), .Y(_15159_) );
	NAND3X1 NAND3X1_3230 ( .gnd(gnd), .vdd(vdd), .A(_15151_), .B(_15150_), .C(_15157_), .Y(_15160_) );
	OAI21X1 OAI21X1_3230 ( .gnd(gnd), .vdd(vdd), .A(_15149_), .B(_15156_), .C(_15153_), .Y(_15161_) );
	AOI21X1 AOI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .B(_15161_), .C(_14834_), .Y(_15162_) );
	NAND2X1 NAND2X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_14842_), .B(_14840_), .Y(_15163_) );
	OAI21X1 OAI21X1_3231 ( .gnd(gnd), .vdd(vdd), .A(_14835_), .B(_14836_), .C(_15163_), .Y(_15164_) );
	OAI21X1 OAI21X1_3232 ( .gnd(gnd), .vdd(vdd), .A(_15159_), .B(_15162_), .C(_15164_), .Y(_15165_) );
	NAND3X1 NAND3X1_3231 ( .gnd(gnd), .vdd(vdd), .A(_14834_), .B(_15161_), .C(_15160_), .Y(_15167_) );
	NOR3X1 NOR3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_15149_), .B(_15153_), .C(_15156_), .Y(_15168_) );
	AOI21X1 AOI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_15150_), .B(_15151_), .C(_15157_), .Y(_15169_) );
	OAI21X1 OAI21X1_3233 ( .gnd(gnd), .vdd(vdd), .A(_15169_), .B(_15168_), .C(_14833_), .Y(_15170_) );
	AOI21X1 AOI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_14842_), .B(_14840_), .C(_14838_), .Y(_15171_) );
	NAND3X1 NAND3X1_3232 ( .gnd(gnd), .vdd(vdd), .A(_15167_), .B(_15171_), .C(_15170_), .Y(_15172_) );
	OAI21X1 OAI21X1_3234 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .B(_14929_), .C(_14926_), .Y(_15173_) );
	NAND3X1 NAND3X1_3233 ( .gnd(gnd), .vdd(vdd), .A(_15165_), .B(_15172_), .C(_15173_), .Y(_15174_) );
	NAND2X1 NAND2X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_15165_), .Y(_15175_) );
	NAND3X1 NAND3X1_3234 ( .gnd(gnd), .vdd(vdd), .A(_14926_), .B(_15175_), .C(_15076_), .Y(_15176_) );
	NAND3X1 NAND3X1_3235 ( .gnd(gnd), .vdd(vdd), .A(_15134_), .B(_15174_), .C(_15176_), .Y(_15178_) );
	INVX1 INVX1_1999 ( .gnd(gnd), .vdd(vdd), .A(_15134_), .Y(_15179_) );
	OR2X2 OR2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .B(_15173_), .Y(_15180_) );
	NAND2X1 NAND2X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_15173_), .B(_15175_), .Y(_15181_) );
	NAND3X1 NAND3X1_3236 ( .gnd(gnd), .vdd(vdd), .A(_15179_), .B(_15181_), .C(_15180_), .Y(_15182_) );
	AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_15182_), .B(_15178_), .Y(_15183_) );
	AOI21X1 AOI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_15063_), .B(_15067_), .C(_14933_), .Y(_15184_) );
	OAI21X1 OAI21X1_3235 ( .gnd(gnd), .vdd(vdd), .A(_15184_), .B(_15078_), .C(_15069_), .Y(_15185_) );
	NAND2X1 NAND2X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_14911_), .B(_14917_), .Y(_15186_) );
	NAND2X1 NAND2X1_3010 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf4), .B(adder_bOperand_23_), .Y(_15187_) );
	INVX1 INVX1_2000 ( .gnd(gnd), .vdd(vdd), .A(_15187_), .Y(_15189_) );
	NAND2X1 NAND2X1_3011 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf0), .B(adder_bOperand_22_bF_buf2), .Y(_15190_) );
	OAI21X1 OAI21X1_3236 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_14862_), .C(_14861_), .Y(_15191_) );
	OAI21X1 OAI21X1_3237 ( .gnd(gnd), .vdd(vdd), .A(_15141_), .B(_15190_), .C(_15191_), .Y(_15192_) );
	XNOR2X1 XNOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_15192_), .B(_15189_), .Y(_15193_) );
	INVX1 INVX1_2001 ( .gnd(gnd), .vdd(vdd), .A(_15193_), .Y(_15194_) );
	NOR2X1 NOR2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_14578_), .B(_14874_), .Y(_15195_) );
	AOI21X1 AOI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_14875_), .B(_14871_), .C(_15195_), .Y(_15196_) );
	INVX1 INVX1_2002 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .Y(_15197_) );
	NAND2X1 NAND2X1_3012 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf3), .B(adder_bOperand_20_bF_buf1), .Y(_15198_) );
	NAND2X1 NAND2X1_3013 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf4), .B(adder_bOperand_19_bF_buf2), .Y(_15200_) );
	OAI21X1 OAI21X1_3238 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_13338_), .C(_14873_), .Y(_15201_) );
	OAI21X1 OAI21X1_3239 ( .gnd(gnd), .vdd(vdd), .A(_14874_), .B(_15200_), .C(_15201_), .Y(_15202_) );
	XOR2X1 XOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_15202_), .B(_15198_), .Y(_15203_) );
	NOR2X1 NOR2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_15197_), .B(_15203_), .Y(_15204_) );
	XNOR2X1 XNOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_15202_), .B(_15198_), .Y(_15205_) );
	NOR2X1 NOR2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .B(_15205_), .Y(_15206_) );
	OAI21X1 OAI21X1_3240 ( .gnd(gnd), .vdd(vdd), .A(_15206_), .B(_15204_), .C(_15194_), .Y(_15207_) );
	NAND2X1 NAND2X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .B(_15205_), .Y(_15208_) );
	NAND2X1 NAND2X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_15197_), .B(_15203_), .Y(_15209_) );
	NAND3X1 NAND3X1_3237 ( .gnd(gnd), .vdd(vdd), .A(_15193_), .B(_15208_), .C(_15209_), .Y(_15211_) );
	AND2X2 AND2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_15207_), .B(_15211_), .Y(_15212_) );
	NOR2X1 NOR2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .B(_14897_), .Y(_15213_) );
	OAI21X1 OAI21X1_3241 ( .gnd(gnd), .vdd(vdd), .A(_14907_), .B(_15213_), .C(_14900_), .Y(_15214_) );
	NAND2X1 NAND2X1_3016 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf1), .B(adder_bOperand_15_bF_buf0), .Y(_15215_) );
	OR2X2 OR2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_14599_), .B(_15215_), .Y(_15216_) );
	OAI21X1 OAI21X1_3242 ( .gnd(gnd), .vdd(vdd), .A(_14893_), .B(_14896_), .C(_15216_), .Y(_15217_) );
	NAND2X1 NAND2X1_3017 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf4), .B(adder_bOperand_17_bF_buf1), .Y(_15218_) );
	NAND2X1 NAND2X1_3018 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf0), .B(adder_bOperand_16_bF_buf0), .Y(_15219_) );
	OAI21X1 OAI21X1_3243 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_12131_), .C(_14894_), .Y(_15220_) );
	OAI21X1 OAI21X1_3244 ( .gnd(gnd), .vdd(vdd), .A(_15215_), .B(_15219_), .C(_15220_), .Y(_15222_) );
	XOR2X1 XOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_15222_), .B(_15218_), .Y(_15223_) );
	OAI21X1 OAI21X1_3245 ( .gnd(gnd), .vdd(vdd), .A(_14960_), .B(_14941_), .C(_14939_), .Y(_15224_) );
	NAND2X1 NAND2X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_15224_), .B(_15223_), .Y(_15225_) );
	AND2X2 AND2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_15222_), .B(_15218_), .Y(_15226_) );
	NOR2X1 NOR2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_15218_), .B(_15222_), .Y(_15227_) );
	INVX1 INVX1_2003 ( .gnd(gnd), .vdd(vdd), .A(_14939_), .Y(_15228_) );
	AOI21X1 AOI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_14935_), .C(_15228_), .Y(_15229_) );
	OAI21X1 OAI21X1_3246 ( .gnd(gnd), .vdd(vdd), .A(_15227_), .B(_15226_), .C(_15229_), .Y(_15230_) );
	NAND3X1 NAND3X1_3238 ( .gnd(gnd), .vdd(vdd), .A(_15217_), .B(_15230_), .C(_15225_), .Y(_15231_) );
	INVX1 INVX1_2004 ( .gnd(gnd), .vdd(vdd), .A(_15217_), .Y(_15233_) );
	NAND2X1 NAND2X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_15229_), .B(_15223_), .Y(_15234_) );
	OAI21X1 OAI21X1_3247 ( .gnd(gnd), .vdd(vdd), .A(_15227_), .B(_15226_), .C(_15224_), .Y(_15235_) );
	NAND3X1 NAND3X1_3239 ( .gnd(gnd), .vdd(vdd), .A(_15233_), .B(_15234_), .C(_15235_), .Y(_15236_) );
	NAND3X1 NAND3X1_3240 ( .gnd(gnd), .vdd(vdd), .A(_15231_), .B(_15236_), .C(_15214_), .Y(_15237_) );
	NOR2X1 NOR2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_14898_), .B(_14904_), .Y(_15238_) );
	AOI21X1 AOI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_14891_), .B(_14905_), .C(_15238_), .Y(_15239_) );
	AOI21X1 AOI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_15235_), .B(_15234_), .C(_15233_), .Y(_15240_) );
	AOI21X1 AOI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_15225_), .B(_15230_), .C(_15217_), .Y(_15241_) );
	OAI21X1 OAI21X1_3248 ( .gnd(gnd), .vdd(vdd), .A(_15241_), .B(_15240_), .C(_15239_), .Y(_15242_) );
	NAND3X1 NAND3X1_3241 ( .gnd(gnd), .vdd(vdd), .A(_15237_), .B(_15242_), .C(_15212_), .Y(_15244_) );
	NAND2X1 NAND2X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_15211_), .B(_15207_), .Y(_15245_) );
	OAI21X1 OAI21X1_3249 ( .gnd(gnd), .vdd(vdd), .A(_15241_), .B(_15240_), .C(_15214_), .Y(_15246_) );
	NAND3X1 NAND3X1_3242 ( .gnd(gnd), .vdd(vdd), .A(_15231_), .B(_15236_), .C(_15239_), .Y(_15247_) );
	NAND3X1 NAND3X1_3243 ( .gnd(gnd), .vdd(vdd), .A(_15245_), .B(_15246_), .C(_15247_), .Y(_15248_) );
	NAND2X1 NAND2X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .B(_14974_), .Y(_15249_) );
	AOI21X1 AOI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_15244_), .B(_15248_), .C(_15249_), .Y(_15250_) );
	NAND2X1 NAND2X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_15248_), .B(_15244_), .Y(_15251_) );
	INVX1 INVX1_2005 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .Y(_15252_) );
	AOI21X1 AOI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_14934_), .B(_14973_), .C(_15252_), .Y(_15253_) );
	NOR2X1 NOR2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_15253_), .B(_15251_), .Y(_15254_) );
	OAI21X1 OAI21X1_3250 ( .gnd(gnd), .vdd(vdd), .A(_15250_), .B(_15254_), .C(_15186_), .Y(_15255_) );
	INVX1 INVX1_2006 ( .gnd(gnd), .vdd(vdd), .A(_15186_), .Y(_15256_) );
	AOI21X1 AOI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_15247_), .B(_15246_), .C(_15245_), .Y(_15257_) );
	AOI21X1 AOI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_15242_), .B(_15237_), .C(_15212_), .Y(_15258_) );
	OAI21X1 OAI21X1_3251 ( .gnd(gnd), .vdd(vdd), .A(_15258_), .B(_15257_), .C(_15253_), .Y(_15259_) );
	NAND3X1 NAND3X1_3244 ( .gnd(gnd), .vdd(vdd), .A(_15248_), .B(_15244_), .C(_15249_), .Y(_15260_) );
	NAND3X1 NAND3X1_3245 ( .gnd(gnd), .vdd(vdd), .A(_15259_), .B(_15256_), .C(_15260_), .Y(_15261_) );
	NAND2X1 NAND2X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_15261_), .B(_15255_), .Y(_15262_) );
	OAI21X1 OAI21X1_3252 ( .gnd(gnd), .vdd(vdd), .A(_15064_), .B(_15065_), .C(_15062_), .Y(_15263_) );
	NAND2X1 NAND2X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14959_), .Y(_15266_) );
	INVX1 INVX1_2007 ( .gnd(gnd), .vdd(vdd), .A(_15266_), .Y(_15267_) );
	NAND2X1 NAND2X1_3026 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf1), .B(aOperand_frameOut_14_bF_buf3), .Y(_15268_) );
	OAI22X1 OAI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(_17157_), .B(_12039_), .C(_11858_), .D(_17319_), .Y(_15269_) );
	OAI21X1 OAI21X1_3253 ( .gnd(gnd), .vdd(vdd), .A(_14937_), .B(_15268_), .C(_15269_), .Y(_15270_) );
	OAI21X1 OAI21X1_3254 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf1), .B(_12365_), .C(_15270_), .Y(_15271_) );
	NAND2X1 NAND2X1_3027 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf4), .B(adder_bOperand_14_bF_buf1), .Y(_15272_) );
	OR2X2 OR2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_15270_), .B(_15272_), .Y(_15273_) );
	NAND2X1 NAND2X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_15271_), .B(_15273_), .Y(_15274_) );
	INVX1 INVX1_2008 ( .gnd(gnd), .vdd(vdd), .A(_15274_), .Y(_15275_) );
	NOR2X1 NOR2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_14654_), .B(_14950_), .Y(_15277_) );
	NAND2X1 NAND2X1_3029 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf2), .B(aOperand_frameOut_15_bF_buf0), .Y(_15278_) );
	NAND2X1 NAND2X1_3030 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf4), .B(aOperand_frameOut_17_bF_buf3), .Y(_15279_) );
	OAI21X1 OAI21X1_3255 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf2), .B(_12708_), .C(_14949_), .Y(_15280_) );
	OAI21X1 OAI21X1_3256 ( .gnd(gnd), .vdd(vdd), .A(_14950_), .B(_15279_), .C(_15280_), .Y(_15281_) );
	XOR2X1 XOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_15281_), .B(_15278_), .Y(_15282_) );
	OAI21X1 OAI21X1_3257 ( .gnd(gnd), .vdd(vdd), .A(_15277_), .B(_14955_), .C(_15282_), .Y(_15283_) );
	NOR2X1 NOR2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_15277_), .B(_14955_), .Y(_15284_) );
	OAI21X1 OAI21X1_3258 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf2), .B(_12233_), .C(_15281_), .Y(_15285_) );
	OR2X2 OR2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_15281_), .B(_15278_), .Y(_15286_) );
	NAND2X1 NAND2X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_15285_), .B(_15286_), .Y(_15288_) );
	NAND2X1 NAND2X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_15284_), .B(_15288_), .Y(_15289_) );
	NAND3X1 NAND3X1_3246 ( .gnd(gnd), .vdd(vdd), .A(_15283_), .B(_15275_), .C(_15289_), .Y(_15290_) );
	OAI21X1 OAI21X1_3259 ( .gnd(gnd), .vdd(vdd), .A(_15277_), .B(_14955_), .C(_15288_), .Y(_15291_) );
	NAND2X1 NAND2X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_15282_), .B(_15284_), .Y(_15292_) );
	NAND3X1 NAND3X1_3247 ( .gnd(gnd), .vdd(vdd), .A(_15274_), .B(_15292_), .C(_15291_), .Y(_15293_) );
	NAND2X1 NAND2X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_15001_), .Y(_15294_) );
	NAND3X1 NAND3X1_3248 ( .gnd(gnd), .vdd(vdd), .A(_15290_), .B(_15293_), .C(_15294_), .Y(_15295_) );
	AOI21X1 AOI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_15291_), .B(_15292_), .C(_15274_), .Y(_15296_) );
	AOI21X1 AOI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_15289_), .B(_15283_), .C(_15275_), .Y(_15297_) );
	AND2X2 AND2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_15001_), .B(_14996_), .Y(_15299_) );
	OAI21X1 OAI21X1_3260 ( .gnd(gnd), .vdd(vdd), .A(_15297_), .B(_15296_), .C(_15299_), .Y(_15300_) );
	NAND3X1 NAND3X1_3249 ( .gnd(gnd), .vdd(vdd), .A(_15267_), .B(_15295_), .C(_15300_), .Y(_15301_) );
	NAND3X1 NAND3X1_3250 ( .gnd(gnd), .vdd(vdd), .A(_15290_), .B(_15293_), .C(_15299_), .Y(_15302_) );
	OAI21X1 OAI21X1_3261 ( .gnd(gnd), .vdd(vdd), .A(_15297_), .B(_15296_), .C(_15294_), .Y(_15303_) );
	NAND3X1 NAND3X1_3251 ( .gnd(gnd), .vdd(vdd), .A(_15266_), .B(_15302_), .C(_15303_), .Y(_15304_) );
	NAND2X1 NAND2X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_15301_), .B(_15304_), .Y(_15305_) );
	OAI21X1 OAI21X1_3262 ( .gnd(gnd), .vdd(vdd), .A(_15059_), .B(_15058_), .C(_15051_), .Y(_15306_) );
	OAI21X1 OAI21X1_3263 ( .gnd(gnd), .vdd(vdd), .A(_14998_), .B(_14985_), .C(_14989_), .Y(_15307_) );
	NAND2X1 NAND2X1_3036 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf1), .B(aOperand_frameOut_18_bF_buf1), .Y(_15308_) );
	NAND2X1 NAND2X1_3037 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf4), .B(aOperand_frameOut_19_bF_buf3), .Y(_15310_) );
	NAND2X1 NAND2X1_3038 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf3), .B(aOperand_frameOut_20_bF_buf0), .Y(_15311_) );
	OAI21X1 OAI21X1_3264 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf1), .B(_13514_), .C(_14984_), .Y(_15312_) );
	OAI21X1 OAI21X1_3265 ( .gnd(gnd), .vdd(vdd), .A(_15310_), .B(_15311_), .C(_15312_), .Y(_15313_) );
	XOR2X1 XOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_15313_), .B(_15308_), .Y(_15314_) );
	NOR2X1 NOR2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_14709_), .B(_15014_), .Y(_15315_) );
	AOI21X1 AOI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_15015_), .B(_15010_), .C(_15315_), .Y(_15316_) );
	INVX1 INVX1_2009 ( .gnd(gnd), .vdd(vdd), .A(_15316_), .Y(_15317_) );
	NAND2X1 NAND2X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_15317_), .B(_15314_), .Y(_15318_) );
	OAI21X1 OAI21X1_3266 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf0), .B(_13796_), .C(_15313_), .Y(_15319_) );
	OR2X2 OR2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_15313_), .B(_15308_), .Y(_15321_) );
	NAND2X1 NAND2X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_15319_), .B(_15321_), .Y(_15322_) );
	NAND2X1 NAND2X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_15316_), .B(_15322_), .Y(_15323_) );
	NAND3X1 NAND3X1_3252 ( .gnd(gnd), .vdd(vdd), .A(_15307_), .B(_15318_), .C(_15323_), .Y(_15324_) );
	INVX1 INVX1_2010 ( .gnd(gnd), .vdd(vdd), .A(_15307_), .Y(_15325_) );
	NAND2X1 NAND2X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_15316_), .B(_15314_), .Y(_15326_) );
	NAND2X1 NAND2X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_15317_), .B(_15322_), .Y(_15327_) );
	NAND3X1 NAND3X1_3253 ( .gnd(gnd), .vdd(vdd), .A(_15325_), .B(_15326_), .C(_15327_), .Y(_15328_) );
	AND2X2 AND2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_15324_), .B(_15328_), .Y(_15329_) );
	NAND2X1 NAND2X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .B(_15049_), .Y(_15330_) );
	NAND2X1 NAND2X1_3045 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf1), .B(aOperand_frameOut_23_), .Y(_15332_) );
	OAI21X1 OAI21X1_3267 ( .gnd(gnd), .vdd(vdd), .A(_11971__bF_buf2), .B(_14436_), .C(_15012_), .Y(_15333_) );
	OAI21X1 OAI21X1_3268 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .B(_15332_), .C(_15333_), .Y(_15334_) );
	OAI21X1 OAI21X1_3269 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf2), .B(_13812_), .C(_15334_), .Y(_15335_) );
	NOR2X1 NOR2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf1), .B(_13812_), .Y(_15336_) );
	INVX1 INVX1_2011 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .Y(_15337_) );
	INVX1 INVX1_2012 ( .gnd(gnd), .vdd(vdd), .A(_15332_), .Y(_15338_) );
	NAND2X1 NAND2X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_15337_), .B(_15338_), .Y(_15339_) );
	NAND3X1 NAND3X1_3254 ( .gnd(gnd), .vdd(vdd), .A(_15336_), .B(_15333_), .C(_15339_), .Y(_15340_) );
	NAND2X1 NAND2X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_15340_), .B(_15335_), .Y(_15341_) );
	INVX1 INVX1_2013 ( .gnd(gnd), .vdd(vdd), .A(_15341_), .Y(_15343_) );
	AOI22X1 AOI22X1_361 ( .gnd(gnd), .vdd(vdd), .A(_15031_), .B(_15032_), .C(_15022_), .D(_15028_), .Y(_15344_) );
	INVX1 INVX1_2014 ( .gnd(gnd), .vdd(vdd), .A(_15344_), .Y(_15345_) );
	NOR2X1 NOR2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_14722_), .Y(_15346_) );
	NAND2X1 NAND2X1_3048 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf6), .B(aOperand_frameOut_25_bF_buf1), .Y(_15347_) );
	NAND2X1 NAND2X1_3049 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf1), .B(aOperand_frameOut_26_), .Y(_15348_) );
	NAND2X1 NAND2X1_3050 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf5), .B(aOperand_frameOut_26_), .Y(_15349_) );
	OAI21X1 OAI21X1_3270 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf3), .B(_15027_), .C(_15349_), .Y(_15350_) );
	OAI21X1 OAI21X1_3271 ( .gnd(gnd), .vdd(vdd), .A(_15347_), .B(_15348_), .C(_15350_), .Y(_15351_) );
	XNOR2X1 XNOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_15351_), .B(_15346_), .Y(_15352_) );
	NAND2X1 NAND2X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_15345_), .B(_15352_), .Y(_15354_) );
	INVX1 INVX1_2015 ( .gnd(gnd), .vdd(vdd), .A(_15346_), .Y(_15355_) );
	NOR2X1 NOR2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_15355_), .B(_15351_), .Y(_15356_) );
	NOR2X1 NOR2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_15026_), .B(_15349_), .Y(_15357_) );
	INVX1 INVX1_2016 ( .gnd(gnd), .vdd(vdd), .A(_15357_), .Y(_15358_) );
	AOI21X1 AOI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_15358_), .B(_15350_), .C(_15346_), .Y(_15359_) );
	OAI21X1 OAI21X1_3272 ( .gnd(gnd), .vdd(vdd), .A(_15356_), .B(_15359_), .C(_15344_), .Y(_15360_) );
	NAND3X1 NAND3X1_3255 ( .gnd(gnd), .vdd(vdd), .A(_15343_), .B(_15360_), .C(_15354_), .Y(_15361_) );
	NOR3X1 NOR3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_15344_), .B(_15356_), .C(_15359_), .Y(_15362_) );
	INVX1 INVX1_2017 ( .gnd(gnd), .vdd(vdd), .A(_15360_), .Y(_15363_) );
	OAI21X1 OAI21X1_3273 ( .gnd(gnd), .vdd(vdd), .A(_15362_), .B(_15363_), .C(_15341_), .Y(_15365_) );
	NAND3X1 NAND3X1_3256 ( .gnd(gnd), .vdd(vdd), .A(_15361_), .B(_15330_), .C(_15365_), .Y(_15366_) );
	INVX1 INVX1_2018 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .Y(_15367_) );
	AOI21X1 AOI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_15041_), .B(_15043_), .C(_15367_), .Y(_15368_) );
	OAI21X1 OAI21X1_3274 ( .gnd(gnd), .vdd(vdd), .A(_15356_), .B(_15359_), .C(_15345_), .Y(_15369_) );
	NAND2X1 NAND2X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_15344_), .B(_15352_), .Y(_15370_) );
	AOI21X1 AOI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_15370_), .B(_15369_), .C(_15341_), .Y(_15371_) );
	AOI21X1 AOI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_15354_), .B(_15360_), .C(_15343_), .Y(_15372_) );
	OAI21X1 OAI21X1_3275 ( .gnd(gnd), .vdd(vdd), .A(_15371_), .B(_15372_), .C(_15368_), .Y(_15373_) );
	NAND3X1 NAND3X1_3257 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15329_), .C(_15373_), .Y(_15374_) );
	NAND2X1 NAND2X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_15328_), .B(_15324_), .Y(_15376_) );
	OAI21X1 OAI21X1_3276 ( .gnd(gnd), .vdd(vdd), .A(_15371_), .B(_15372_), .C(_15330_), .Y(_15377_) );
	NAND3X1 NAND3X1_3258 ( .gnd(gnd), .vdd(vdd), .A(_15368_), .B(_15361_), .C(_15365_), .Y(_15378_) );
	NAND3X1 NAND3X1_3259 ( .gnd(gnd), .vdd(vdd), .A(_15376_), .B(_15378_), .C(_15377_), .Y(_15379_) );
	NAND3X1 NAND3X1_3260 ( .gnd(gnd), .vdd(vdd), .A(_15379_), .B(_15374_), .C(_15306_), .Y(_15380_) );
	AOI21X1 AOI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .B(_15045_), .C(_15060_), .Y(_15381_) );
	AOI21X1 AOI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_15377_), .B(_15378_), .C(_15376_), .Y(_15382_) );
	AOI21X1 AOI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_15373_), .B(_15366_), .C(_15329_), .Y(_15383_) );
	OAI21X1 OAI21X1_3277 ( .gnd(gnd), .vdd(vdd), .A(_15382_), .B(_15383_), .C(_15381_), .Y(_15384_) );
	NAND3X1 NAND3X1_3261 ( .gnd(gnd), .vdd(vdd), .A(_15305_), .B(_15380_), .C(_15384_), .Y(_15385_) );
	AND2X2 AND2X2_378 ( .gnd(gnd), .vdd(vdd), .A(_15304_), .B(_15301_), .Y(_15387_) );
	OAI21X1 OAI21X1_3278 ( .gnd(gnd), .vdd(vdd), .A(_15382_), .B(_15383_), .C(_15306_), .Y(_15388_) );
	NAND3X1 NAND3X1_3262 ( .gnd(gnd), .vdd(vdd), .A(_15381_), .B(_15379_), .C(_15374_), .Y(_15389_) );
	NAND3X1 NAND3X1_3263 ( .gnd(gnd), .vdd(vdd), .A(_15389_), .B(_15388_), .C(_15387_), .Y(_15390_) );
	NAND3X1 NAND3X1_3264 ( .gnd(gnd), .vdd(vdd), .A(_15385_), .B(_15263_), .C(_15390_), .Y(_15391_) );
	AOI21X1 AOI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_14979_), .B(_15055_), .C(_15066_), .Y(_15392_) );
	AOI21X1 AOI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_15388_), .B(_15389_), .C(_15387_), .Y(_15393_) );
	AOI21X1 AOI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_15384_), .B(_15380_), .C(_15305_), .Y(_15394_) );
	OAI21X1 OAI21X1_3279 ( .gnd(gnd), .vdd(vdd), .A(_15393_), .B(_15394_), .C(_15392_), .Y(_15395_) );
	NAND3X1 NAND3X1_3265 ( .gnd(gnd), .vdd(vdd), .A(_15391_), .B(_15395_), .C(_15262_), .Y(_15396_) );
	NAND3X1 NAND3X1_3266 ( .gnd(gnd), .vdd(vdd), .A(_15186_), .B(_15259_), .C(_15260_), .Y(_15398_) );
	OAI21X1 OAI21X1_3280 ( .gnd(gnd), .vdd(vdd), .A(_15250_), .B(_15254_), .C(_15256_), .Y(_15399_) );
	NAND2X1 NAND2X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_15398_), .B(_15399_), .Y(_15400_) );
	OAI21X1 OAI21X1_3281 ( .gnd(gnd), .vdd(vdd), .A(_15393_), .B(_15394_), .C(_15263_), .Y(_15401_) );
	NAND3X1 NAND3X1_3267 ( .gnd(gnd), .vdd(vdd), .A(_15385_), .B(_15390_), .C(_15392_), .Y(_15402_) );
	NAND3X1 NAND3X1_3268 ( .gnd(gnd), .vdd(vdd), .A(_15402_), .B(_15401_), .C(_15400_), .Y(_15403_) );
	NAND3X1 NAND3X1_3269 ( .gnd(gnd), .vdd(vdd), .A(_15396_), .B(_15403_), .C(_15185_), .Y(_15404_) );
	NOR3X1 NOR3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_15071_), .B(_15073_), .C(_15072_), .Y(_15405_) );
	AOI21X1 AOI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .B(_14932_), .C(_15405_), .Y(_15406_) );
	AOI21X1 AOI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_15401_), .B(_15402_), .C(_15400_), .Y(_15407_) );
	AOI21X1 AOI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_15395_), .B(_15391_), .C(_15262_), .Y(_15409_) );
	OAI21X1 OAI21X1_3282 ( .gnd(gnd), .vdd(vdd), .A(_15407_), .B(_15409_), .C(_15406_), .Y(_15410_) );
	NAND3X1 NAND3X1_3270 ( .gnd(gnd), .vdd(vdd), .A(_15404_), .B(_15410_), .C(_15183_), .Y(_15411_) );
	NAND2X1 NAND2X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_15178_), .B(_15182_), .Y(_15412_) );
	OAI21X1 OAI21X1_3283 ( .gnd(gnd), .vdd(vdd), .A(_15407_), .B(_15409_), .C(_15185_), .Y(_15413_) );
	NAND3X1 NAND3X1_3271 ( .gnd(gnd), .vdd(vdd), .A(_15396_), .B(_15403_), .C(_15406_), .Y(_15414_) );
	NAND3X1 NAND3X1_3272 ( .gnd(gnd), .vdd(vdd), .A(_15412_), .B(_15414_), .C(_15413_), .Y(_15415_) );
	NAND3X1 NAND3X1_3273 ( .gnd(gnd), .vdd(vdd), .A(_15415_), .B(_15411_), .C(_15132_), .Y(_15416_) );
	NOR3X1 NOR3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_15085_), .B(_15086_), .C(_15087_), .Y(_15417_) );
	AOI21X1 AOI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_14854_), .B(_15088_), .C(_15417_), .Y(_15418_) );
	AOI21X1 AOI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_15413_), .B(_15414_), .C(_15412_), .Y(_15420_) );
	AOI21X1 AOI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_15410_), .B(_15404_), .C(_15183_), .Y(_15421_) );
	OAI21X1 OAI21X1_3284 ( .gnd(gnd), .vdd(vdd), .A(_15420_), .B(_15421_), .C(_15418_), .Y(_15422_) );
	NAND3X1 NAND3X1_3274 ( .gnd(gnd), .vdd(vdd), .A(_15130_), .B(_15416_), .C(_15422_), .Y(_15423_) );
	INVX1 INVX1_2019 ( .gnd(gnd), .vdd(vdd), .A(_15130_), .Y(_15424_) );
	OAI21X1 OAI21X1_3285 ( .gnd(gnd), .vdd(vdd), .A(_15420_), .B(_15421_), .C(_15132_), .Y(_15425_) );
	NAND3X1 NAND3X1_3275 ( .gnd(gnd), .vdd(vdd), .A(_15411_), .B(_15415_), .C(_15418_), .Y(_15426_) );
	NAND3X1 NAND3X1_3276 ( .gnd(gnd), .vdd(vdd), .A(_15424_), .B(_15425_), .C(_15426_), .Y(_15427_) );
	NAND3X1 NAND3X1_3277 ( .gnd(gnd), .vdd(vdd), .A(_15423_), .B(_15129_), .C(_15427_), .Y(_15428_) );
	INVX1 INVX1_2020 ( .gnd(gnd), .vdd(vdd), .A(_15097_), .Y(_15429_) );
	AOI21X1 AOI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_14817_), .B(_15103_), .C(_15429_), .Y(_15431_) );
	AOI21X1 AOI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_15426_), .B(_15425_), .C(_15424_), .Y(_15432_) );
	AOI21X1 AOI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_15422_), .B(_15416_), .C(_15130_), .Y(_15433_) );
	OAI21X1 OAI21X1_3286 ( .gnd(gnd), .vdd(vdd), .A(_15433_), .B(_15432_), .C(_15431_), .Y(_15434_) );
	NAND3X1 NAND3X1_3278 ( .gnd(gnd), .vdd(vdd), .A(_15108_), .B(_15428_), .C(_15434_), .Y(_15435_) );
	NOR3X1 NOR3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_15110_), .B(_15113_), .C(_15111_), .Y(_15436_) );
	OAI21X1 OAI21X1_3287 ( .gnd(gnd), .vdd(vdd), .A(_15433_), .B(_15432_), .C(_15129_), .Y(_15437_) );
	NAND3X1 NAND3X1_3279 ( .gnd(gnd), .vdd(vdd), .A(_15423_), .B(_15427_), .C(_15431_), .Y(_15438_) );
	NAND3X1 NAND3X1_3280 ( .gnd(gnd), .vdd(vdd), .A(_15437_), .B(_15438_), .C(_15436_), .Y(_15439_) );
	NAND2X1 NAND2X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_15435_), .B(_15439_), .Y(_15440_) );
	XOR2X1 XOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_15127_), .B(_15440_), .Y(mulOut_26_) );
	AOI21X1 AOI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_15438_), .B(_15437_), .C(_15108_), .Y(_15442_) );
	INVX1 INVX1_2021 ( .gnd(gnd), .vdd(vdd), .A(_15442_), .Y(_15443_) );
	NOR2X1 NOR2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_15113_), .B(_15111_), .Y(_15444_) );
	AOI22X1 AOI22X1_362 ( .gnd(gnd), .vdd(vdd), .A(_15444_), .B(_14816_), .C(_15437_), .D(_15438_), .Y(_15445_) );
	AOI21X1 AOI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_15434_), .B(_15428_), .C(_15108_), .Y(_15446_) );
	OAI21X1 OAI21X1_3288 ( .gnd(gnd), .vdd(vdd), .A(_15445_), .B(_15446_), .C(_15127_), .Y(_15447_) );
	AOI21X1 AOI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_15411_), .B(_15415_), .C(_15132_), .Y(_15448_) );
	OAI21X1 OAI21X1_3289 ( .gnd(gnd), .vdd(vdd), .A(_15424_), .B(_15448_), .C(_15416_), .Y(_15449_) );
	NAND2X1 NAND2X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15178_), .Y(_15450_) );
	AOI21X1 AOI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_15396_), .B(_15403_), .C(_15185_), .Y(_15452_) );
	OAI21X1 OAI21X1_3290 ( .gnd(gnd), .vdd(vdd), .A(_15412_), .B(_15452_), .C(_15404_), .Y(_15453_) );
	INVX1 INVX1_2022 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_27_), .Y(_15454_) );
	NOR2X1 NOR2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf1), .B(_15454_), .Y(_15455_) );
	AOI21X1 AOI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14834_), .C(_15168_), .Y(_15456_) );
	OAI21X1 OAI21X1_3291 ( .gnd(gnd), .vdd(vdd), .A(_15147_), .B(_15143_), .C(_15151_), .Y(_15457_) );
	NAND2X1 NAND2X1_3058 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf2), .B(adder_bOperand_24_), .Y(_15458_) );
	NOR2X1 NOR2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_14823_), .B(_15458_), .Y(_15459_) );
	NOR2X1 NOR2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_15136_), .B(_15139_), .Y(_15460_) );
	NOR2X1 NOR2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_15459_), .B(_15460_), .Y(_15461_) );
	NAND2X1 NAND2X1_3059 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf3), .B(adder_bOperand_26_), .Y(_15463_) );
	OAI21X1 OAI21X1_3292 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_14544_), .C(_15137_), .Y(_15464_) );
	NAND2X1 NAND2X1_3060 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf3), .B(adder_bOperand_25_), .Y(_15465_) );
	OAI21X1 OAI21X1_3293 ( .gnd(gnd), .vdd(vdd), .A(_15458_), .B(_15465_), .C(_15464_), .Y(_15466_) );
	XOR2X1 XOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_15466_), .B(_15463_), .Y(_15467_) );
	OAI22X1 OAI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_15141_), .B(_15190_), .C(_15187_), .D(_15192_), .Y(_15468_) );
	INVX1 INVX1_2023 ( .gnd(gnd), .vdd(vdd), .A(_15468_), .Y(_15469_) );
	NAND2X1 NAND2X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_15467_), .B(_15469_), .Y(_15470_) );
	AND2X2 AND2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_15466_), .B(_15463_), .Y(_15471_) );
	NOR2X1 NOR2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_15463_), .B(_15466_), .Y(_15472_) );
	OAI21X1 OAI21X1_3294 ( .gnd(gnd), .vdd(vdd), .A(_15472_), .B(_15471_), .C(_15468_), .Y(_15474_) );
	AOI21X1 AOI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_15470_), .B(_15474_), .C(_15461_), .Y(_15475_) );
	INVX1 INVX1_2024 ( .gnd(gnd), .vdd(vdd), .A(_15461_), .Y(_15476_) );
	NAND2X1 NAND2X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_15468_), .B(_15467_), .Y(_15477_) );
	OAI21X1 OAI21X1_3295 ( .gnd(gnd), .vdd(vdd), .A(_15472_), .B(_15471_), .C(_15469_), .Y(_15478_) );
	AOI21X1 AOI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_15478_), .B(_15477_), .C(_15476_), .Y(_15479_) );
	AOI21X1 AOI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_15193_), .B(_15208_), .C(_15206_), .Y(_15480_) );
	OAI21X1 OAI21X1_3296 ( .gnd(gnd), .vdd(vdd), .A(_15475_), .B(_15479_), .C(_15480_), .Y(_15481_) );
	NAND3X1 NAND3X1_3281 ( .gnd(gnd), .vdd(vdd), .A(_15477_), .B(_15476_), .C(_15478_), .Y(_15482_) );
	NAND3X1 NAND3X1_3282 ( .gnd(gnd), .vdd(vdd), .A(_15461_), .B(_15474_), .C(_15470_), .Y(_15483_) );
	OAI21X1 OAI21X1_3297 ( .gnd(gnd), .vdd(vdd), .A(_15194_), .B(_15204_), .C(_15209_), .Y(_15485_) );
	NAND3X1 NAND3X1_3283 ( .gnd(gnd), .vdd(vdd), .A(_15482_), .B(_15483_), .C(_15485_), .Y(_15486_) );
	AOI21X1 AOI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_15481_), .B(_15486_), .C(_15457_), .Y(_15487_) );
	NAND3X1 NAND3X1_3284 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .B(_15486_), .C(_15481_), .Y(_15488_) );
	INVX1 INVX1_2025 ( .gnd(gnd), .vdd(vdd), .A(_15488_), .Y(_15489_) );
	OAI21X1 OAI21X1_3298 ( .gnd(gnd), .vdd(vdd), .A(_15487_), .B(_15489_), .C(_15456_), .Y(_15490_) );
	OAI21X1 OAI21X1_3299 ( .gnd(gnd), .vdd(vdd), .A(_14833_), .B(_15169_), .C(_15160_), .Y(_15491_) );
	INVX1 INVX1_2026 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .Y(_15492_) );
	AOI21X1 AOI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_15482_), .B(_15483_), .C(_15485_), .Y(_15493_) );
	INVX1 INVX1_2027 ( .gnd(gnd), .vdd(vdd), .A(_15486_), .Y(_15494_) );
	OAI21X1 OAI21X1_3300 ( .gnd(gnd), .vdd(vdd), .A(_15493_), .B(_15494_), .C(_15492_), .Y(_15496_) );
	NAND3X1 NAND3X1_3285 ( .gnd(gnd), .vdd(vdd), .A(_15488_), .B(_15496_), .C(_15491_), .Y(_15497_) );
	AOI21X1 AOI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_15490_), .B(_15497_), .C(_15455_), .Y(_15498_) );
	INVX1 INVX1_2028 ( .gnd(gnd), .vdd(vdd), .A(_15498_), .Y(_15499_) );
	NAND3X1 NAND3X1_3286 ( .gnd(gnd), .vdd(vdd), .A(_15455_), .B(_15497_), .C(_15490_), .Y(_15500_) );
	OAI21X1 OAI21X1_3301 ( .gnd(gnd), .vdd(vdd), .A(_15256_), .B(_15250_), .C(_15260_), .Y(_15501_) );
	NAND3X1 NAND3X1_3287 ( .gnd(gnd), .vdd(vdd), .A(_15500_), .B(_15501_), .C(_15499_), .Y(_15502_) );
	INVX1 INVX1_2029 ( .gnd(gnd), .vdd(vdd), .A(_15500_), .Y(_15503_) );
	INVX1 INVX1_2030 ( .gnd(gnd), .vdd(vdd), .A(_15501_), .Y(_15504_) );
	OAI21X1 OAI21X1_3302 ( .gnd(gnd), .vdd(vdd), .A(_15498_), .B(_15503_), .C(_15504_), .Y(_15505_) );
	NAND3X1 NAND3X1_3288 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_15502_), .C(_15505_), .Y(_15507_) );
	INVX1 INVX1_2031 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .Y(_15508_) );
	OAI21X1 OAI21X1_3303 ( .gnd(gnd), .vdd(vdd), .A(_15498_), .B(_15503_), .C(_15501_), .Y(_15509_) );
	NAND3X1 NAND3X1_3289 ( .gnd(gnd), .vdd(vdd), .A(_15500_), .B(_15504_), .C(_15499_), .Y(_15510_) );
	NAND3X1 NAND3X1_3290 ( .gnd(gnd), .vdd(vdd), .A(_15508_), .B(_15510_), .C(_15509_), .Y(_15511_) );
	NAND2X1 NAND2X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_15507_), .B(_15511_), .Y(_15512_) );
	AOI21X1 AOI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_15390_), .B(_15385_), .C(_15263_), .Y(_15513_) );
	OAI21X1 OAI21X1_3304 ( .gnd(gnd), .vdd(vdd), .A(_15513_), .B(_15400_), .C(_15391_), .Y(_15514_) );
	NAND2X1 NAND2X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_15237_), .B(_15244_), .Y(_15515_) );
	INVX1 INVX1_2032 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .Y(_15516_) );
	NOR2X1 NOR2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf2), .B(_14564_), .Y(_15518_) );
	NAND2X1 NAND2X1_3065 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf2), .B(adder_bOperand_21_bF_buf1), .Y(_15519_) );
	NOR2X1 NOR2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_15190_), .B(_15519_), .Y(_15520_) );
	AND2X2 AND2X2_380 ( .gnd(gnd), .vdd(vdd), .A(_15190_), .B(_15519_), .Y(_15521_) );
	NOR2X1 NOR2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_15520_), .B(_15521_), .Y(_15522_) );
	OR2X2 OR2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_15522_), .B(_15518_), .Y(_15523_) );
	NAND2X1 NAND2X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_15518_), .B(_15522_), .Y(_15524_) );
	NAND2X1 NAND2X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_15524_), .B(_15523_), .Y(_15525_) );
	INVX1 INVX1_2033 ( .gnd(gnd), .vdd(vdd), .A(_15525_), .Y(_15526_) );
	NOR2X1 NOR2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_14874_), .B(_15200_), .Y(_15527_) );
	NOR2X1 NOR2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_15198_), .B(_15202_), .Y(_15529_) );
	OR2X2 OR2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_15529_), .B(_15527_), .Y(_15530_) );
	NAND2X1 NAND2X1_3068 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf3), .B(adder_bOperand_18_bF_buf2), .Y(_15531_) );
	XNOR2X1 XNOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .B(_15531_), .Y(_15532_) );
	OAI21X1 OAI21X1_3305 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_13334_), .C(_15532_), .Y(_15533_) );
	NAND2X1 NAND2X1_3069 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf4), .B(adder_bOperand_20_bF_buf0), .Y(_15534_) );
	OR2X2 OR2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_15532_), .B(_15534_), .Y(_15535_) );
	NAND3X1 NAND3X1_3291 ( .gnd(gnd), .vdd(vdd), .A(_15533_), .B(_15535_), .C(_15530_), .Y(_15536_) );
	NOR2X1 NOR2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_15527_), .B(_15529_), .Y(_15537_) );
	NAND2X1 NAND2X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_15533_), .B(_15535_), .Y(_15538_) );
	NAND2X1 NAND2X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_15537_), .B(_15538_), .Y(_15540_) );
	NAND3X1 NAND3X1_3292 ( .gnd(gnd), .vdd(vdd), .A(_15526_), .B(_15540_), .C(_15536_), .Y(_15541_) );
	NAND2X1 NAND2X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_15540_), .B(_15536_), .Y(_15542_) );
	NAND2X1 NAND2X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_15525_), .B(_15542_), .Y(_15543_) );
	AND2X2 AND2X2_381 ( .gnd(gnd), .vdd(vdd), .A(_15543_), .B(_15541_), .Y(_15544_) );
	NAND2X1 NAND2X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_15225_), .B(_15231_), .Y(_15545_) );
	NAND2X1 NAND2X1_3075 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf4), .B(adder_bOperand_15_bF_buf4), .Y(_15546_) );
	OR2X2 OR2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .B(_15546_), .Y(_15547_) );
	OAI21X1 OAI21X1_3306 ( .gnd(gnd), .vdd(vdd), .A(_15218_), .B(_15222_), .C(_15547_), .Y(_15548_) );
	OAI21X1 OAI21X1_3307 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf0), .B(_12131_), .C(_15219_), .Y(_15549_) );
	NAND2X1 NAND2X1_3076 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf3), .B(adder_bOperand_16_bF_buf3), .Y(_15550_) );
	OAI21X1 OAI21X1_3308 ( .gnd(gnd), .vdd(vdd), .A(_15546_), .B(_15550_), .C(_15549_), .Y(_15551_) );
	OAI21X1 OAI21X1_3309 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_12566_), .C(_15551_), .Y(_15552_) );
	NAND2X1 NAND2X1_3077 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf0), .B(adder_bOperand_17_bF_buf0), .Y(_15553_) );
	OR2X2 OR2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_15551_), .B(_15553_), .Y(_15554_) );
	AND2X2 AND2X2_382 ( .gnd(gnd), .vdd(vdd), .A(_15554_), .B(_15552_), .Y(_15555_) );
	OR2X2 OR2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_14937_), .B(_15268_), .Y(_15556_) );
	OAI21X1 OAI21X1_3310 ( .gnd(gnd), .vdd(vdd), .A(_15272_), .B(_15270_), .C(_15556_), .Y(_15557_) );
	NAND2X1 NAND2X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_15557_), .B(_15555_), .Y(_15558_) );
	NAND2X1 NAND2X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_15552_), .B(_15554_), .Y(_15559_) );
	INVX1 INVX1_2034 ( .gnd(gnd), .vdd(vdd), .A(_15557_), .Y(_15561_) );
	NAND2X1 NAND2X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_15561_), .B(_15559_), .Y(_15562_) );
	NAND3X1 NAND3X1_3293 ( .gnd(gnd), .vdd(vdd), .A(_15548_), .B(_15562_), .C(_15558_), .Y(_15563_) );
	INVX1 INVX1_2035 ( .gnd(gnd), .vdd(vdd), .A(_15548_), .Y(_15564_) );
	NAND2X1 NAND2X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_15562_), .B(_15558_), .Y(_15565_) );
	NAND2X1 NAND2X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_15564_), .B(_15565_), .Y(_15566_) );
	NAND3X1 NAND3X1_3294 ( .gnd(gnd), .vdd(vdd), .A(_15545_), .B(_15563_), .C(_15566_), .Y(_15567_) );
	AND2X2 AND2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_15231_), .B(_15225_), .Y(_15568_) );
	NAND2X1 NAND2X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_15561_), .B(_15555_), .Y(_15569_) );
	NAND2X1 NAND2X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_15557_), .B(_15559_), .Y(_15570_) );
	AOI21X1 AOI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_15569_), .B(_15570_), .C(_15564_), .Y(_15573_) );
	AOI21X1 AOI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_15558_), .B(_15562_), .C(_15548_), .Y(_15574_) );
	OAI21X1 OAI21X1_3311 ( .gnd(gnd), .vdd(vdd), .A(_15573_), .B(_15574_), .C(_15568_), .Y(_15575_) );
	NAND3X1 NAND3X1_3295 ( .gnd(gnd), .vdd(vdd), .A(_15575_), .B(_15567_), .C(_15544_), .Y(_15576_) );
	NAND2X1 NAND2X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_15541_), .B(_15543_), .Y(_15577_) );
	OAI21X1 OAI21X1_3312 ( .gnd(gnd), .vdd(vdd), .A(_15573_), .B(_15574_), .C(_15545_), .Y(_15578_) );
	NAND3X1 NAND3X1_3296 ( .gnd(gnd), .vdd(vdd), .A(_15563_), .B(_15568_), .C(_15566_), .Y(_15579_) );
	NAND3X1 NAND3X1_3297 ( .gnd(gnd), .vdd(vdd), .A(_15578_), .B(_15577_), .C(_15579_), .Y(_15580_) );
	NAND3X1 NAND3X1_3298 ( .gnd(gnd), .vdd(vdd), .A(_15266_), .B(_15295_), .C(_15300_), .Y(_15581_) );
	NAND2X1 NAND2X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_15295_), .B(_15581_), .Y(_15582_) );
	NAND3X1 NAND3X1_3299 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .B(_15576_), .C(_15582_), .Y(_15584_) );
	AOI21X1 AOI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_15579_), .B(_15578_), .C(_15577_), .Y(_15585_) );
	AOI21X1 AOI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_15567_), .B(_15575_), .C(_15544_), .Y(_15586_) );
	AND2X2 AND2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_15581_), .B(_15295_), .Y(_15587_) );
	OAI21X1 OAI21X1_3313 ( .gnd(gnd), .vdd(vdd), .A(_15585_), .B(_15586_), .C(_15587_), .Y(_15588_) );
	NAND3X1 NAND3X1_3300 ( .gnd(gnd), .vdd(vdd), .A(_15516_), .B(_15584_), .C(_15588_), .Y(_15589_) );
	NAND3X1 NAND3X1_3301 ( .gnd(gnd), .vdd(vdd), .A(_15576_), .B(_15580_), .C(_15587_), .Y(_15590_) );
	OAI21X1 OAI21X1_3314 ( .gnd(gnd), .vdd(vdd), .A(_15585_), .B(_15586_), .C(_15582_), .Y(_15591_) );
	NAND3X1 NAND3X1_3302 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .B(_15591_), .C(_15590_), .Y(_15592_) );
	NAND2X1 NAND2X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_15589_), .B(_15592_), .Y(_15593_) );
	AOI21X1 AOI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_15374_), .B(_15379_), .C(_15306_), .Y(_15595_) );
	OAI21X1 OAI21X1_3315 ( .gnd(gnd), .vdd(vdd), .A(_15595_), .B(_15387_), .C(_15380_), .Y(_15596_) );
	OAI21X1 OAI21X1_3316 ( .gnd(gnd), .vdd(vdd), .A(_15284_), .B(_15288_), .C(_15290_), .Y(_15597_) );
	INVX1 INVX1_2036 ( .gnd(gnd), .vdd(vdd), .A(_15597_), .Y(_15598_) );
	NOR2X1 NOR2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_11858_), .B(_12365_), .Y(_15599_) );
	NAND2X1 NAND2X1_3088 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf0), .B(aOperand_frameOut_15_bF_buf4), .Y(_15600_) );
	AND2X2 AND2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_15268_), .B(_15600_), .Y(_15601_) );
	NOR2X1 NOR2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_15268_), .B(_15600_), .Y(_15602_) );
	NOR2X1 NOR2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_15602_), .B(_15601_), .Y(_15603_) );
	OR2X2 OR2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_15603_), .B(_15599_), .Y(_15604_) );
	NAND2X1 NAND2X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_15599_), .B(_15603_), .Y(_15606_) );
	NAND2X1 NAND2X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_15606_), .B(_15604_), .Y(_15607_) );
	INVX1 INVX1_2037 ( .gnd(gnd), .vdd(vdd), .A(_15607_), .Y(_15608_) );
	NAND2X1 NAND2X1_3091 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf1), .B(aOperand_frameOut_17_bF_buf2), .Y(_15609_) );
	OR2X2 OR2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_14949_), .B(_15609_), .Y(_15610_) );
	OAI21X1 OAI21X1_3317 ( .gnd(gnd), .vdd(vdd), .A(_15278_), .B(_15281_), .C(_15610_), .Y(_15611_) );
	OAI21X1 OAI21X1_3318 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf1), .B(_13796_), .C(_15279_), .Y(_15612_) );
	NAND2X1 NAND2X1_3092 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf3), .B(aOperand_frameOut_18_bF_buf0), .Y(_15613_) );
	OAI21X1 OAI21X1_3319 ( .gnd(gnd), .vdd(vdd), .A(_15609_), .B(_15613_), .C(_15612_), .Y(_15614_) );
	OAI21X1 OAI21X1_3320 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf1), .B(_12461_), .C(_15614_), .Y(_15615_) );
	NAND2X1 NAND2X1_3093 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf1), .B(aOperand_frameOut_16_bF_buf3), .Y(_15617_) );
	OR2X2 OR2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_15614_), .B(_15617_), .Y(_15618_) );
	AND2X2 AND2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_15618_), .B(_15615_), .Y(_15619_) );
	NAND2X1 NAND2X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_15611_), .B(_15619_), .Y(_15620_) );
	INVX1 INVX1_2038 ( .gnd(gnd), .vdd(vdd), .A(_15611_), .Y(_15621_) );
	NAND2X1 NAND2X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_15615_), .B(_15618_), .Y(_15622_) );
	NAND2X1 NAND2X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_15621_), .B(_15622_), .Y(_15623_) );
	NAND3X1 NAND3X1_3303 ( .gnd(gnd), .vdd(vdd), .A(_15623_), .B(_15608_), .C(_15620_), .Y(_15624_) );
	NAND2X1 NAND2X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_15623_), .B(_15620_), .Y(_15625_) );
	NAND2X1 NAND2X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_15607_), .B(_15625_), .Y(_15626_) );
	OAI21X1 OAI21X1_3321 ( .gnd(gnd), .vdd(vdd), .A(_15322_), .B(_15316_), .C(_15324_), .Y(_15628_) );
	NAND3X1 NAND3X1_3304 ( .gnd(gnd), .vdd(vdd), .A(_15624_), .B(_15628_), .C(_15626_), .Y(_15629_) );
	INVX1 INVX1_2039 ( .gnd(gnd), .vdd(vdd), .A(_15624_), .Y(_15630_) );
	AOI21X1 AOI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_15620_), .B(_15623_), .C(_15608_), .Y(_15631_) );
	AND2X2 AND2X2_387 ( .gnd(gnd), .vdd(vdd), .A(_15324_), .B(_15318_), .Y(_15632_) );
	OAI21X1 OAI21X1_3322 ( .gnd(gnd), .vdd(vdd), .A(_15631_), .B(_15630_), .C(_15632_), .Y(_15633_) );
	NAND3X1 NAND3X1_3305 ( .gnd(gnd), .vdd(vdd), .A(_15598_), .B(_15629_), .C(_15633_), .Y(_15634_) );
	NAND3X1 NAND3X1_3306 ( .gnd(gnd), .vdd(vdd), .A(_15624_), .B(_15626_), .C(_15632_), .Y(_15635_) );
	OAI21X1 OAI21X1_3323 ( .gnd(gnd), .vdd(vdd), .A(_15631_), .B(_15630_), .C(_15628_), .Y(_15636_) );
	NAND3X1 NAND3X1_3307 ( .gnd(gnd), .vdd(vdd), .A(_15597_), .B(_15635_), .C(_15636_), .Y(_15637_) );
	NAND2X1 NAND2X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_15634_), .B(_15637_), .Y(_15639_) );
	AOI21X1 AOI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_15365_), .B(_15361_), .C(_15330_), .Y(_15640_) );
	OAI21X1 OAI21X1_3324 ( .gnd(gnd), .vdd(vdd), .A(_15376_), .B(_15640_), .C(_15366_), .Y(_15641_) );
	NAND2X1 NAND2X1_3100 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf3), .B(aOperand_frameOut_20_bF_buf4), .Y(_15642_) );
	OR2X2 OR2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .B(_15642_), .Y(_15643_) );
	OAI21X1 OAI21X1_3325 ( .gnd(gnd), .vdd(vdd), .A(_15308_), .B(_15313_), .C(_15643_), .Y(_15644_) );
	INVX1 INVX1_2040 ( .gnd(gnd), .vdd(vdd), .A(_15644_), .Y(_15645_) );
	NAND2X1 NAND2X1_3101 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf0), .B(aOperand_frameOut_19_bF_buf2), .Y(_15646_) );
	OAI21X1 OAI21X1_3326 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf0), .B(_13812_), .C(_15311_), .Y(_15647_) );
	NAND2X1 NAND2X1_3102 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf2), .B(aOperand_frameOut_21_bF_buf3), .Y(_15648_) );
	OAI21X1 OAI21X1_3327 ( .gnd(gnd), .vdd(vdd), .A(_15642_), .B(_15648_), .C(_15647_), .Y(_15649_) );
	XOR2X1 XOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_15649_), .B(_15646_), .Y(_15650_) );
	OAI21X1 OAI21X1_3328 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .B(_15332_), .C(_15340_), .Y(_15651_) );
	NOR2X1 NOR2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_15651_), .B(_15650_), .Y(_15652_) );
	AND2X2 AND2X2_388 ( .gnd(gnd), .vdd(vdd), .A(_15650_), .B(_15651_), .Y(_15653_) );
	OAI21X1 OAI21X1_3329 ( .gnd(gnd), .vdd(vdd), .A(_15652_), .B(_15653_), .C(_15645_), .Y(_15654_) );
	OR2X2 OR2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_15650_), .B(_15651_), .Y(_15655_) );
	NAND2X1 NAND2X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_15651_), .B(_15650_), .Y(_15656_) );
	NAND3X1 NAND3X1_3308 ( .gnd(gnd), .vdd(vdd), .A(_15644_), .B(_15656_), .C(_15655_), .Y(_15657_) );
	NAND2X1 NAND2X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_15657_), .B(_15654_), .Y(_15658_) );
	OAI21X1 OAI21X1_3330 ( .gnd(gnd), .vdd(vdd), .A(_15341_), .B(_15363_), .C(_15354_), .Y(_15660_) );
	NOR2X1 NOR2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf0), .B(_14125_), .Y(_15661_) );
	INVX1 INVX1_2041 ( .gnd(gnd), .vdd(vdd), .A(_15661_), .Y(_15662_) );
	NAND2X1 NAND2X1_3105 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf1), .B(aOperand_frameOut_24_bF_buf3), .Y(_15663_) );
	AND2X2 AND2X2_389 ( .gnd(gnd), .vdd(vdd), .A(_15332_), .B(_15663_), .Y(_15664_) );
	NOR2X1 NOR2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_15332_), .B(_15663_), .Y(_15665_) );
	OAI21X1 OAI21X1_3331 ( .gnd(gnd), .vdd(vdd), .A(_15665_), .B(_15664_), .C(_15662_), .Y(_15666_) );
	NOR2X1 NOR2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_15665_), .B(_15664_), .Y(_15667_) );
	NAND2X1 NAND2X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_15661_), .B(_15667_), .Y(_15668_) );
	NAND2X1 NAND2X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_15666_), .B(_15668_), .Y(_15669_) );
	AOI21X1 AOI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_15350_), .B(_15346_), .C(_15357_), .Y(_15671_) );
	INVX1 INVX1_2042 ( .gnd(gnd), .vdd(vdd), .A(_15671_), .Y(_15672_) );
	NAND2X1 NAND2X1_3108 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf0), .B(aOperand_frameOut_27_), .Y(_15673_) );
	INVX1 INVX1_2043 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_26_), .Y(_15674_) );
	NAND2X1 NAND2X1_3109 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf4), .B(aOperand_frameOut_27_), .Y(_15675_) );
	OAI21X1 OAI21X1_3332 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf2), .B(_15674_), .C(_15675_), .Y(_15676_) );
	OAI21X1 OAI21X1_3333 ( .gnd(gnd), .vdd(vdd), .A(_15349_), .B(_15673_), .C(_15676_), .Y(_15677_) );
	OAI21X1 OAI21X1_3334 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_15027_), .C(_15677_), .Y(_15678_) );
	NAND2X1 NAND2X1_3110 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf1), .B(aOperand_frameOut_25_bF_buf0), .Y(_15679_) );
	OR2X2 OR2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_15677_), .B(_15679_), .Y(_15680_) );
	AOI21X1 AOI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_15680_), .B(_15678_), .C(_15672_), .Y(_15682_) );
	AND2X2 AND2X2_390 ( .gnd(gnd), .vdd(vdd), .A(_15677_), .B(_15679_), .Y(_15683_) );
	NOR2X1 NOR2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_15679_), .B(_15677_), .Y(_15684_) );
	NOR3X1 NOR3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_15671_), .B(_15684_), .C(_15683_), .Y(_15685_) );
	OAI21X1 OAI21X1_3335 ( .gnd(gnd), .vdd(vdd), .A(_15682_), .B(_15685_), .C(_15669_), .Y(_15686_) );
	INVX1 INVX1_2044 ( .gnd(gnd), .vdd(vdd), .A(_15669_), .Y(_15687_) );
	OAI21X1 OAI21X1_3336 ( .gnd(gnd), .vdd(vdd), .A(_15684_), .B(_15683_), .C(_15671_), .Y(_15688_) );
	NAND3X1 NAND3X1_3309 ( .gnd(gnd), .vdd(vdd), .A(_15678_), .B(_15672_), .C(_15680_), .Y(_15689_) );
	NAND3X1 NAND3X1_3310 ( .gnd(gnd), .vdd(vdd), .A(_15688_), .B(_15689_), .C(_15687_), .Y(_15690_) );
	AOI21X1 AOI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_15686_), .B(_15690_), .C(_15660_), .Y(_15691_) );
	AOI21X1 AOI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_15343_), .B(_15360_), .C(_15362_), .Y(_15693_) );
	AOI21X1 AOI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_15688_), .B(_15689_), .C(_15687_), .Y(_15694_) );
	NOR3X1 NOR3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_15669_), .B(_15682_), .C(_15685_), .Y(_15695_) );
	NOR3X1 NOR3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_15693_), .B(_15694_), .C(_15695_), .Y(_15696_) );
	OAI21X1 OAI21X1_3337 ( .gnd(gnd), .vdd(vdd), .A(_15691_), .B(_15696_), .C(_15658_), .Y(_15697_) );
	AND2X2 AND2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_15654_), .B(_15657_), .Y(_15698_) );
	OAI21X1 OAI21X1_3338 ( .gnd(gnd), .vdd(vdd), .A(_15694_), .B(_15695_), .C(_15693_), .Y(_15699_) );
	NAND3X1 NAND3X1_3311 ( .gnd(gnd), .vdd(vdd), .A(_15686_), .B(_15690_), .C(_15660_), .Y(_15700_) );
	NAND3X1 NAND3X1_3312 ( .gnd(gnd), .vdd(vdd), .A(_15700_), .B(_15699_), .C(_15698_), .Y(_15701_) );
	NAND3X1 NAND3X1_3313 ( .gnd(gnd), .vdd(vdd), .A(_15701_), .B(_15641_), .C(_15697_), .Y(_15702_) );
	INVX1 INVX1_2045 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .Y(_15704_) );
	AOI21X1 AOI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_15329_), .B(_15373_), .C(_15704_), .Y(_15705_) );
	AOI21X1 AOI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_15699_), .B(_15700_), .C(_15698_), .Y(_15706_) );
	NOR3X1 NOR3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_15658_), .B(_15691_), .C(_15696_), .Y(_15707_) );
	OAI21X1 OAI21X1_3339 ( .gnd(gnd), .vdd(vdd), .A(_15706_), .B(_15707_), .C(_15705_), .Y(_15708_) );
	NAND3X1 NAND3X1_3314 ( .gnd(gnd), .vdd(vdd), .A(_15702_), .B(_15708_), .C(_15639_), .Y(_15709_) );
	NAND3X1 NAND3X1_3315 ( .gnd(gnd), .vdd(vdd), .A(_15597_), .B(_15629_), .C(_15633_), .Y(_15710_) );
	NAND3X1 NAND3X1_3316 ( .gnd(gnd), .vdd(vdd), .A(_15598_), .B(_15635_), .C(_15636_), .Y(_15711_) );
	NAND2X1 NAND2X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_15710_), .B(_15711_), .Y(_15712_) );
	OAI21X1 OAI21X1_3340 ( .gnd(gnd), .vdd(vdd), .A(_15706_), .B(_15707_), .C(_15641_), .Y(_15713_) );
	NAND3X1 NAND3X1_3317 ( .gnd(gnd), .vdd(vdd), .A(_15697_), .B(_15701_), .C(_15705_), .Y(_15715_) );
	NAND3X1 NAND3X1_3318 ( .gnd(gnd), .vdd(vdd), .A(_15715_), .B(_15713_), .C(_15712_), .Y(_15716_) );
	NAND3X1 NAND3X1_3319 ( .gnd(gnd), .vdd(vdd), .A(_15596_), .B(_15709_), .C(_15716_), .Y(_15717_) );
	INVX1 INVX1_2046 ( .gnd(gnd), .vdd(vdd), .A(_15380_), .Y(_15718_) );
	AOI21X1 AOI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_15305_), .B(_15384_), .C(_15718_), .Y(_15719_) );
	AOI22X1 AOI22X1_363 ( .gnd(gnd), .vdd(vdd), .A(_15634_), .B(_15637_), .C(_15715_), .D(_15713_), .Y(_15720_) );
	AOI22X1 AOI22X1_364 ( .gnd(gnd), .vdd(vdd), .A(_15710_), .B(_15711_), .C(_15702_), .D(_15708_), .Y(_15721_) );
	OAI21X1 OAI21X1_3341 ( .gnd(gnd), .vdd(vdd), .A(_15720_), .B(_15721_), .C(_15719_), .Y(_15722_) );
	NAND3X1 NAND3X1_3320 ( .gnd(gnd), .vdd(vdd), .A(_15717_), .B(_15722_), .C(_15593_), .Y(_15723_) );
	NAND3X1 NAND3X1_3321 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .B(_15584_), .C(_15588_), .Y(_15724_) );
	NAND3X1 NAND3X1_3322 ( .gnd(gnd), .vdd(vdd), .A(_15516_), .B(_15591_), .C(_15590_), .Y(_15726_) );
	NAND2X1 NAND2X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_15724_), .B(_15726_), .Y(_15727_) );
	OAI21X1 OAI21X1_3342 ( .gnd(gnd), .vdd(vdd), .A(_15720_), .B(_15721_), .C(_15596_), .Y(_15728_) );
	NAND3X1 NAND3X1_3323 ( .gnd(gnd), .vdd(vdd), .A(_15719_), .B(_15709_), .C(_15716_), .Y(_15729_) );
	NAND3X1 NAND3X1_3324 ( .gnd(gnd), .vdd(vdd), .A(_15729_), .B(_15728_), .C(_15727_), .Y(_15730_) );
	NAND3X1 NAND3X1_3325 ( .gnd(gnd), .vdd(vdd), .A(_15514_), .B(_15723_), .C(_15730_), .Y(_15731_) );
	INVX1 INVX1_2047 ( .gnd(gnd), .vdd(vdd), .A(_15391_), .Y(_15732_) );
	AOI21X1 AOI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_15262_), .B(_15395_), .C(_15732_), .Y(_15733_) );
	AOI22X1 AOI22X1_365 ( .gnd(gnd), .vdd(vdd), .A(_15589_), .B(_15592_), .C(_15729_), .D(_15728_), .Y(_15734_) );
	AOI22X1 AOI22X1_366 ( .gnd(gnd), .vdd(vdd), .A(_15724_), .B(_15726_), .C(_15717_), .D(_15722_), .Y(_15735_) );
	OAI21X1 OAI21X1_3343 ( .gnd(gnd), .vdd(vdd), .A(_15734_), .B(_15735_), .C(_15733_), .Y(_15737_) );
	NAND3X1 NAND3X1_3326 ( .gnd(gnd), .vdd(vdd), .A(_15731_), .B(_15737_), .C(_15512_), .Y(_15738_) );
	NAND3X1 NAND3X1_3327 ( .gnd(gnd), .vdd(vdd), .A(_15508_), .B(_15502_), .C(_15505_), .Y(_15739_) );
	NAND3X1 NAND3X1_3328 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_15510_), .C(_15509_), .Y(_15740_) );
	NAND2X1 NAND2X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_15739_), .B(_15740_), .Y(_15741_) );
	OAI21X1 OAI21X1_3344 ( .gnd(gnd), .vdd(vdd), .A(_15734_), .B(_15735_), .C(_15514_), .Y(_15742_) );
	NAND3X1 NAND3X1_3329 ( .gnd(gnd), .vdd(vdd), .A(_15723_), .B(_15730_), .C(_15733_), .Y(_15743_) );
	NAND3X1 NAND3X1_3330 ( .gnd(gnd), .vdd(vdd), .A(_15743_), .B(_15742_), .C(_15741_), .Y(_15744_) );
	NAND3X1 NAND3X1_3331 ( .gnd(gnd), .vdd(vdd), .A(_15453_), .B(_15738_), .C(_15744_), .Y(_15745_) );
	INVX1 INVX1_2048 ( .gnd(gnd), .vdd(vdd), .A(_15404_), .Y(_15746_) );
	AOI21X1 AOI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .B(_15410_), .C(_15746_), .Y(_15748_) );
	AOI22X1 AOI22X1_367 ( .gnd(gnd), .vdd(vdd), .A(_15507_), .B(_15511_), .C(_15743_), .D(_15742_), .Y(_15749_) );
	AOI22X1 AOI22X1_368 ( .gnd(gnd), .vdd(vdd), .A(_15739_), .B(_15740_), .C(_15731_), .D(_15737_), .Y(_15750_) );
	OAI21X1 OAI21X1_3345 ( .gnd(gnd), .vdd(vdd), .A(_15749_), .B(_15750_), .C(_15748_), .Y(_15751_) );
	NAND3X1 NAND3X1_3332 ( .gnd(gnd), .vdd(vdd), .A(_15450_), .B(_15745_), .C(_15751_), .Y(_15752_) );
	INVX1 INVX1_2049 ( .gnd(gnd), .vdd(vdd), .A(_15450_), .Y(_15753_) );
	OAI21X1 OAI21X1_3346 ( .gnd(gnd), .vdd(vdd), .A(_15749_), .B(_15750_), .C(_15453_), .Y(_15754_) );
	NAND3X1 NAND3X1_3333 ( .gnd(gnd), .vdd(vdd), .A(_15738_), .B(_15744_), .C(_15748_), .Y(_15755_) );
	NAND3X1 NAND3X1_3334 ( .gnd(gnd), .vdd(vdd), .A(_15753_), .B(_15755_), .C(_15754_), .Y(_15756_) );
	NAND3X1 NAND3X1_3335 ( .gnd(gnd), .vdd(vdd), .A(_15449_), .B(_15752_), .C(_15756_), .Y(_15757_) );
	INVX1 INVX1_2050 ( .gnd(gnd), .vdd(vdd), .A(_15416_), .Y(_15759_) );
	AOI21X1 AOI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_15130_), .B(_15422_), .C(_15759_), .Y(_15760_) );
	AOI22X1 AOI22X1_369 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15178_), .C(_15755_), .D(_15754_), .Y(_15761_) );
	AOI21X1 AOI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_15751_), .B(_15745_), .C(_15450_), .Y(_15762_) );
	OAI21X1 OAI21X1_3347 ( .gnd(gnd), .vdd(vdd), .A(_15761_), .B(_15762_), .C(_15760_), .Y(_15763_) );
	NAND3X1 NAND3X1_3336 ( .gnd(gnd), .vdd(vdd), .A(_15428_), .B(_15757_), .C(_15763_), .Y(_15764_) );
	INVX1 INVX1_2051 ( .gnd(gnd), .vdd(vdd), .A(_15428_), .Y(_15765_) );
	OAI21X1 OAI21X1_3348 ( .gnd(gnd), .vdd(vdd), .A(_15761_), .B(_15762_), .C(_15449_), .Y(_15766_) );
	NAND3X1 NAND3X1_3337 ( .gnd(gnd), .vdd(vdd), .A(_15752_), .B(_15756_), .C(_15760_), .Y(_15767_) );
	NAND3X1 NAND3X1_3338 ( .gnd(gnd), .vdd(vdd), .A(_15766_), .B(_15767_), .C(_15765_), .Y(_15768_) );
	NAND2X1 NAND2X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_15764_), .B(_15768_), .Y(_15770_) );
	NAND3X1 NAND3X1_3339 ( .gnd(gnd), .vdd(vdd), .A(_15443_), .B(_15770_), .C(_15447_), .Y(_15771_) );
	AND2X2 AND2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_15127_), .B(_15440_), .Y(_15772_) );
	NAND3X1 NAND3X1_3340 ( .gnd(gnd), .vdd(vdd), .A(_15757_), .B(_15763_), .C(_15765_), .Y(_15773_) );
	NAND3X1 NAND3X1_3341 ( .gnd(gnd), .vdd(vdd), .A(_15428_), .B(_15767_), .C(_15766_), .Y(_15774_) );
	NAND2X1 NAND2X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_15774_), .B(_15773_), .Y(_15775_) );
	OAI21X1 OAI21X1_3349 ( .gnd(gnd), .vdd(vdd), .A(_15442_), .B(_15772_), .C(_15775_), .Y(_15776_) );
	NAND2X1 NAND2X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_15771_), .B(_15776_), .Y(mulOut_27_) );
	AOI22X1 AOI22X1_370 ( .gnd(gnd), .vdd(vdd), .A(_14804_), .B(_14809_), .C(_15115_), .D(_15119_), .Y(_15777_) );
	NAND3X1 NAND3X1_3342 ( .gnd(gnd), .vdd(vdd), .A(_15440_), .B(_15777_), .C(_15770_), .Y(_15778_) );
	NAND2X1 NAND2X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_15121_), .B(_15124_), .Y(_15780_) );
	NOR2X1 NOR2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_15433_), .B(_15432_), .Y(_15781_) );
	AOI22X1 AOI22X1_371 ( .gnd(gnd), .vdd(vdd), .A(_15129_), .B(_15781_), .C(_15767_), .D(_15766_), .Y(_15782_) );
	AOI21X1 AOI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_15763_), .B(_15757_), .C(_15428_), .Y(_15783_) );
	OAI22X1 OAI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(_15446_), .B(_15445_), .C(_15782_), .D(_15783_), .Y(_15784_) );
	INVX1 INVX1_2052 ( .gnd(gnd), .vdd(vdd), .A(_15784_), .Y(_15785_) );
	OAI21X1 OAI21X1_3350 ( .gnd(gnd), .vdd(vdd), .A(_15443_), .B(_15775_), .C(_15773_), .Y(_15786_) );
	AOI21X1 AOI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_15785_), .B(_15780_), .C(_15786_), .Y(_15787_) );
	OAI21X1 OAI21X1_3351 ( .gnd(gnd), .vdd(vdd), .A(_15778_), .B(_14539_), .C(_15787_), .Y(_15788_) );
	INVX1 INVX1_2053 ( .gnd(gnd), .vdd(vdd), .A(_15757_), .Y(_15789_) );
	NAND2X1 NAND2X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_15745_), .B(_15752_), .Y(_15791_) );
	NAND2X1 NAND2X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_15502_), .B(_15739_), .Y(_15792_) );
	NAND2X1 NAND2X1_3120 ( .gnd(gnd), .vdd(vdd), .A(_15731_), .B(_15738_), .Y(_15793_) );
	NAND2X1 NAND2X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_15497_), .B(_15500_), .Y(_15794_) );
	INVX1 INVX1_2054 ( .gnd(gnd), .vdd(vdd), .A(_15794_), .Y(_15795_) );
	INVX1 INVX1_2055 ( .gnd(gnd), .vdd(vdd), .A(_15455_), .Y(_15796_) );
	NAND2X1 NAND2X1_3122 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf2), .B(adder_bOperand_28_), .Y(_15797_) );
	INVX1 INVX1_2056 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_28_), .Y(_15798_) );
	OAI22X1 OAI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(_17306__bF_buf0), .B(_15798_), .C(_11874_), .D(_15454_), .Y(_15799_) );
	OAI21X1 OAI21X1_3352 ( .gnd(gnd), .vdd(vdd), .A(_15797_), .B(_15796_), .C(_15799_), .Y(_15800_) );
	INVX1 INVX1_2057 ( .gnd(gnd), .vdd(vdd), .A(_15800_), .Y(_15802_) );
	OAI21X1 OAI21X1_3353 ( .gnd(gnd), .vdd(vdd), .A(_15493_), .B(_15492_), .C(_15486_), .Y(_15803_) );
	NAND2X1 NAND2X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_15477_), .B(_15482_), .Y(_15804_) );
	OAI22X1 OAI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_15458_), .B(_15465_), .C(_15463_), .D(_15466_), .Y(_15805_) );
	INVX1 INVX1_2058 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_26_), .Y(_15806_) );
	NAND2X1 NAND2X1_3124 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf2), .B(adder_bOperand_24_), .Y(_15807_) );
	NAND2X1 NAND2X1_3125 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf0), .B(adder_bOperand_25_), .Y(_15808_) );
	OAI21X1 OAI21X1_3354 ( .gnd(gnd), .vdd(vdd), .A(_12353__bF_buf1), .B(_14544_), .C(_15465_), .Y(_15809_) );
	OAI21X1 OAI21X1_3355 ( .gnd(gnd), .vdd(vdd), .A(_15807_), .B(_15808_), .C(_15809_), .Y(_15810_) );
	OAI21X1 OAI21X1_3356 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf1), .B(_15806_), .C(_15810_), .Y(_15811_) );
	NAND2X1 NAND2X1_3126 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf1), .B(adder_bOperand_26_), .Y(_15813_) );
	OR2X2 OR2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_15810_), .B(_15813_), .Y(_15814_) );
	OAI21X1 OAI21X1_3357 ( .gnd(gnd), .vdd(vdd), .A(_15190_), .B(_15519_), .C(_15524_), .Y(_15815_) );
	NAND3X1 NAND3X1_3343 ( .gnd(gnd), .vdd(vdd), .A(_15811_), .B(_15814_), .C(_15815_), .Y(_15816_) );
	NAND2X1 NAND2X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_15811_), .B(_15814_), .Y(_15817_) );
	AOI21X1 AOI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_15522_), .B(_15518_), .C(_15520_), .Y(_15818_) );
	NAND2X1 NAND2X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_15818_), .B(_15817_), .Y(_15819_) );
	NAND2X1 NAND2X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_15819_), .B(_15816_), .Y(_15820_) );
	XNOR2X1 XNOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_15820_), .B(_15805_), .Y(_15821_) );
	OAI21X1 OAI21X1_3358 ( .gnd(gnd), .vdd(vdd), .A(_15537_), .B(_15538_), .C(_15541_), .Y(_15822_) );
	XOR2X1 XOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_15821_), .B(_15822_), .Y(_15824_) );
	NAND2X1 NAND2X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_15804_), .B(_15824_), .Y(_15825_) );
	INVX1 INVX1_2059 ( .gnd(gnd), .vdd(vdd), .A(_15804_), .Y(_15826_) );
	NAND2X1 NAND2X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_15822_), .B(_15821_), .Y(_15827_) );
	XOR2X1 XOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_15820_), .B(_15805_), .Y(_15828_) );
	NAND3X1 NAND3X1_3344 ( .gnd(gnd), .vdd(vdd), .A(_15536_), .B(_15541_), .C(_15828_), .Y(_15829_) );
	NAND2X1 NAND2X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_15827_), .B(_15829_), .Y(_15830_) );
	NAND2X1 NAND2X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_15826_), .B(_15830_), .Y(_15831_) );
	NAND3X1 NAND3X1_3345 ( .gnd(gnd), .vdd(vdd), .A(_15803_), .B(_15831_), .C(_15825_), .Y(_15832_) );
	INVX1 INVX1_2060 ( .gnd(gnd), .vdd(vdd), .A(_15803_), .Y(_15833_) );
	NOR2X1 NOR2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_15826_), .B(_15830_), .Y(_15835_) );
	NOR2X1 NOR2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_15804_), .B(_15824_), .Y(_15836_) );
	OAI21X1 OAI21X1_3359 ( .gnd(gnd), .vdd(vdd), .A(_15835_), .B(_15836_), .C(_15833_), .Y(_15837_) );
	NAND3X1 NAND3X1_3346 ( .gnd(gnd), .vdd(vdd), .A(_15802_), .B(_15832_), .C(_15837_), .Y(_15838_) );
	OAI21X1 OAI21X1_3360 ( .gnd(gnd), .vdd(vdd), .A(_15835_), .B(_15836_), .C(_15803_), .Y(_15839_) );
	NAND3X1 NAND3X1_3347 ( .gnd(gnd), .vdd(vdd), .A(_15833_), .B(_15831_), .C(_15825_), .Y(_15840_) );
	NAND3X1 NAND3X1_3348 ( .gnd(gnd), .vdd(vdd), .A(_15800_), .B(_15840_), .C(_15839_), .Y(_15841_) );
	NAND2X1 NAND2X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15724_), .Y(_15842_) );
	NAND3X1 NAND3X1_3349 ( .gnd(gnd), .vdd(vdd), .A(_15842_), .B(_15838_), .C(_15841_), .Y(_15843_) );
	AOI21X1 AOI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_15839_), .B(_15840_), .C(_15800_), .Y(_15844_) );
	AOI21X1 AOI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_15837_), .B(_15832_), .C(_15802_), .Y(_15846_) );
	INVX1 INVX1_2061 ( .gnd(gnd), .vdd(vdd), .A(_15842_), .Y(_15847_) );
	OAI21X1 OAI21X1_3361 ( .gnd(gnd), .vdd(vdd), .A(_15844_), .B(_15846_), .C(_15847_), .Y(_15848_) );
	NAND3X1 NAND3X1_3350 ( .gnd(gnd), .vdd(vdd), .A(_15795_), .B(_15843_), .C(_15848_), .Y(_15849_) );
	NAND3X1 NAND3X1_3351 ( .gnd(gnd), .vdd(vdd), .A(_15838_), .B(_15841_), .C(_15847_), .Y(_15850_) );
	OAI21X1 OAI21X1_3362 ( .gnd(gnd), .vdd(vdd), .A(_15844_), .B(_15846_), .C(_15842_), .Y(_15851_) );
	NAND3X1 NAND3X1_3352 ( .gnd(gnd), .vdd(vdd), .A(_15794_), .B(_15850_), .C(_15851_), .Y(_15852_) );
	NAND2X1 NAND2X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_15849_), .B(_15852_), .Y(_15853_) );
	NAND2X1 NAND2X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_15717_), .B(_15723_), .Y(_15854_) );
	NAND2X1 NAND2X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_15567_), .B(_15576_), .Y(_15855_) );
	NOR2X1 NOR2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_14564_), .Y(_15857_) );
	NAND2X1 NAND2X1_3138 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf1), .B(adder_bOperand_22_bF_buf1), .Y(_15858_) );
	NAND2X1 NAND2X1_3139 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf3), .B(adder_bOperand_21_bF_buf0), .Y(_15859_) );
	XOR2X1 XOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_15858_), .B(_15859_), .Y(_15860_) );
	XOR2X1 XOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_15860_), .B(_15857_), .Y(_15861_) );
	OAI21X1 OAI21X1_3363 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .B(_15531_), .C(_15535_), .Y(_15862_) );
	NAND2X1 NAND2X1_3140 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf4), .B(adder_bOperand_19_bF_buf1), .Y(_15863_) );
	NAND2X1 NAND2X1_3141 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf3), .B(adder_bOperand_18_bF_buf1), .Y(_15864_) );
	OAI21X1 OAI21X1_3364 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf0), .B(_13067_), .C(_15864_), .Y(_15865_) );
	OAI21X1 OAI21X1_3365 ( .gnd(gnd), .vdd(vdd), .A(_15531_), .B(_15863_), .C(_15865_), .Y(_15866_) );
	OAI21X1 OAI21X1_3366 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_13334_), .C(_15866_), .Y(_15868_) );
	NAND2X1 NAND2X1_3142 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf3), .B(adder_bOperand_20_bF_buf3), .Y(_15869_) );
	OR2X2 OR2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_15866_), .B(_15869_), .Y(_15870_) );
	NAND2X1 NAND2X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_15868_), .B(_15870_), .Y(_15871_) );
	XNOR2X1 XNOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_15862_), .B(_15871_), .Y(_15872_) );
	NAND2X1 NAND2X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_15861_), .B(_15872_), .Y(_15873_) );
	OR2X2 OR2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_15872_), .B(_15861_), .Y(_15874_) );
	AND2X2 AND2X2_393 ( .gnd(gnd), .vdd(vdd), .A(_15874_), .B(_15873_), .Y(_15875_) );
	OAI21X1 OAI21X1_3367 ( .gnd(gnd), .vdd(vdd), .A(_15559_), .B(_15561_), .C(_15563_), .Y(_15876_) );
	NAND2X1 NAND2X1_3145 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf2), .B(adder_bOperand_15_bF_buf3), .Y(_15877_) );
	OR2X2 OR2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_15219_), .B(_15877_), .Y(_15879_) );
	OAI21X1 OAI21X1_3368 ( .gnd(gnd), .vdd(vdd), .A(_15553_), .B(_15551_), .C(_15879_), .Y(_15880_) );
	NAND2X1 NAND2X1_3146 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf1), .B(adder_bOperand_16_bF_buf2), .Y(_15881_) );
	OAI21X1 OAI21X1_3369 ( .gnd(gnd), .vdd(vdd), .A(_11858_), .B(_12131_), .C(_15550_), .Y(_15882_) );
	OAI21X1 OAI21X1_3370 ( .gnd(gnd), .vdd(vdd), .A(_15877_), .B(_15881_), .C(_15882_), .Y(_15883_) );
	OAI21X1 OAI21X1_3371 ( .gnd(gnd), .vdd(vdd), .A(_17077_), .B(_12566_), .C(_15883_), .Y(_15884_) );
	NAND2X1 NAND2X1_3147 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf3), .B(adder_bOperand_17_bF_buf3), .Y(_15885_) );
	OR2X2 OR2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_15883_), .B(_15885_), .Y(_15886_) );
	NAND2X1 NAND2X1_3148 ( .gnd(gnd), .vdd(vdd), .A(_15884_), .B(_15886_), .Y(_15887_) );
	AOI21X1 AOI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_15603_), .B(_15599_), .C(_15602_), .Y(_15888_) );
	OR2X2 OR2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_15887_), .B(_15888_), .Y(_15890_) );
	NAND2X1 NAND2X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_15888_), .B(_15887_), .Y(_15891_) );
	NAND2X1 NAND2X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_15891_), .B(_15890_), .Y(_15892_) );
	XNOR2X1 XNOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_15892_), .B(_15880_), .Y(_15893_) );
	NAND2X1 NAND2X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_15876_), .B(_15893_), .Y(_15894_) );
	INVX1 INVX1_2062 ( .gnd(gnd), .vdd(vdd), .A(_15876_), .Y(_15895_) );
	INVX1 INVX1_2063 ( .gnd(gnd), .vdd(vdd), .A(_15880_), .Y(_15896_) );
	XNOR2X1 XNOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_15892_), .B(_15896_), .Y(_15897_) );
	NAND2X1 NAND2X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_15895_), .B(_15897_), .Y(_15898_) );
	NAND3X1 NAND3X1_3353 ( .gnd(gnd), .vdd(vdd), .A(_15875_), .B(_15898_), .C(_15894_), .Y(_15899_) );
	NAND2X1 NAND2X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_15873_), .B(_15874_), .Y(_15901_) );
	NAND2X1 NAND2X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_15876_), .B(_15897_), .Y(_15902_) );
	NAND2X1 NAND2X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_15895_), .B(_15893_), .Y(_15903_) );
	NAND3X1 NAND3X1_3354 ( .gnd(gnd), .vdd(vdd), .A(_15901_), .B(_15902_), .C(_15903_), .Y(_15904_) );
	NAND2X1 NAND2X1_3156 ( .gnd(gnd), .vdd(vdd), .A(_15629_), .B(_15710_), .Y(_15905_) );
	NAND3X1 NAND3X1_3355 ( .gnd(gnd), .vdd(vdd), .A(_15905_), .B(_15899_), .C(_15904_), .Y(_15906_) );
	AOI21X1 AOI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_15903_), .B(_15902_), .C(_15901_), .Y(_15907_) );
	AOI21X1 AOI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_15894_), .B(_15898_), .C(_15875_), .Y(_15908_) );
	AND2X2 AND2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_15710_), .B(_15629_), .Y(_15909_) );
	OAI21X1 OAI21X1_3372 ( .gnd(gnd), .vdd(vdd), .A(_15908_), .B(_15907_), .C(_15909_), .Y(_15910_) );
	NAND3X1 NAND3X1_3356 ( .gnd(gnd), .vdd(vdd), .A(_15855_), .B(_15906_), .C(_15910_), .Y(_15912_) );
	INVX1 INVX1_2064 ( .gnd(gnd), .vdd(vdd), .A(_15855_), .Y(_15913_) );
	NAND3X1 NAND3X1_3357 ( .gnd(gnd), .vdd(vdd), .A(_15899_), .B(_15904_), .C(_15909_), .Y(_15914_) );
	OAI21X1 OAI21X1_3373 ( .gnd(gnd), .vdd(vdd), .A(_15908_), .B(_15907_), .C(_15905_), .Y(_15915_) );
	NAND3X1 NAND3X1_3358 ( .gnd(gnd), .vdd(vdd), .A(_15913_), .B(_15914_), .C(_15915_), .Y(_15916_) );
	AND2X2 AND2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_15916_), .B(_15912_), .Y(_15917_) );
	INVX1 INVX1_2065 ( .gnd(gnd), .vdd(vdd), .A(_15702_), .Y(_15918_) );
	AOI21X1 AOI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_15639_), .B(_15708_), .C(_15918_), .Y(_15919_) );
	OAI21X1 OAI21X1_3374 ( .gnd(gnd), .vdd(vdd), .A(_15621_), .B(_15622_), .C(_15624_), .Y(_15920_) );
	NOR2X1 NOR2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_12039_), .B(_12365_), .Y(_15921_) );
	NAND2X1 NAND2X1_3157 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf0), .B(aOperand_frameOut_15_bF_buf3), .Y(_15923_) );
	NAND2X1 NAND2X1_3158 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf3), .B(aOperand_frameOut_16_bF_buf2), .Y(_15924_) );
	XOR2X1 XOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_15923_), .B(_15924_), .Y(_15925_) );
	XOR2X1 XOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_15925_), .B(_15921_), .Y(_15926_) );
	NAND2X1 NAND2X1_3159 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf0), .B(aOperand_frameOut_18_bF_buf4), .Y(_15927_) );
	NOR2X1 NOR2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_15279_), .B(_15927_), .Y(_15928_) );
	NOR2X1 NOR2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_15617_), .B(_15614_), .Y(_15929_) );
	NAND2X1 NAND2X1_3160 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf0), .B(aOperand_frameOut_17_bF_buf1), .Y(_15930_) );
	NAND2X1 NAND2X1_3161 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf2), .B(aOperand_frameOut_19_bF_buf1), .Y(_15931_) );
	OAI21X1 OAI21X1_3375 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf0), .B(_13224_), .C(_15613_), .Y(_15932_) );
	OAI21X1 OAI21X1_3376 ( .gnd(gnd), .vdd(vdd), .A(_15927_), .B(_15931_), .C(_15932_), .Y(_15934_) );
	XOR2X1 XOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_15934_), .B(_15930_), .Y(_15935_) );
	OAI21X1 OAI21X1_3377 ( .gnd(gnd), .vdd(vdd), .A(_15928_), .B(_15929_), .C(_15935_), .Y(_15936_) );
	NOR2X1 NOR2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_15928_), .B(_15929_), .Y(_15937_) );
	OAI21X1 OAI21X1_3378 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf0), .B(_12708_), .C(_15934_), .Y(_15938_) );
	OR2X2 OR2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_15934_), .B(_15930_), .Y(_15939_) );
	NAND2X1 NAND2X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_15938_), .B(_15939_), .Y(_15940_) );
	NAND2X1 NAND2X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_15937_), .B(_15940_), .Y(_15941_) );
	NAND3X1 NAND3X1_3359 ( .gnd(gnd), .vdd(vdd), .A(_15926_), .B(_15936_), .C(_15941_), .Y(_15942_) );
	INVX1 INVX1_2066 ( .gnd(gnd), .vdd(vdd), .A(_15926_), .Y(_15943_) );
	OAI21X1 OAI21X1_3379 ( .gnd(gnd), .vdd(vdd), .A(_15928_), .B(_15929_), .C(_15940_), .Y(_15945_) );
	NAND2X1 NAND2X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_15935_), .B(_15937_), .Y(_15946_) );
	NAND3X1 NAND3X1_3360 ( .gnd(gnd), .vdd(vdd), .A(_15946_), .B(_15943_), .C(_15945_), .Y(_15947_) );
	NAND2X1 NAND2X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_15942_), .B(_15947_), .Y(_15948_) );
	NAND3X1 NAND3X1_3361 ( .gnd(gnd), .vdd(vdd), .A(_15656_), .B(_15657_), .C(_15948_), .Y(_15949_) );
	OAI21X1 OAI21X1_3380 ( .gnd(gnd), .vdd(vdd), .A(_15645_), .B(_15652_), .C(_15656_), .Y(_15950_) );
	NAND3X1 NAND3X1_3362 ( .gnd(gnd), .vdd(vdd), .A(_15942_), .B(_15947_), .C(_15950_), .Y(_15951_) );
	NAND2X1 NAND2X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_15951_), .B(_15949_), .Y(_15952_) );
	XNOR2X1 XNOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_15952_), .B(_15920_), .Y(_15953_) );
	OAI21X1 OAI21X1_3381 ( .gnd(gnd), .vdd(vdd), .A(_15658_), .B(_15691_), .C(_15700_), .Y(_15954_) );
	INVX1 INVX1_2067 ( .gnd(gnd), .vdd(vdd), .A(_15954_), .Y(_15956_) );
	NAND2X1 NAND2X1_3167 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf2), .B(aOperand_frameOut_21_bF_buf2), .Y(_15957_) );
	NOR2X1 NOR2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_15311_), .B(_15957_), .Y(_15958_) );
	NOR2X1 NOR2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_15646_), .B(_15649_), .Y(_15959_) );
	OR2X2 OR2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_15959_), .B(_15958_), .Y(_15960_) );
	NAND2X1 NAND2X1_3168 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf4), .B(aOperand_frameOut_20_bF_buf3), .Y(_15961_) );
	NAND2X1 NAND2X1_3169 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf1), .B(aOperand_frameOut_22_bF_buf1), .Y(_15962_) );
	OAI21X1 OAI21X1_3382 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf3), .B(_14125_), .C(_15648_), .Y(_15963_) );
	OAI21X1 OAI21X1_3383 ( .gnd(gnd), .vdd(vdd), .A(_15957_), .B(_15962_), .C(_15963_), .Y(_15964_) );
	XNOR2X1 XNOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_15964_), .B(_15961_), .Y(_15965_) );
	AOI21X1 AOI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_15667_), .B(_15661_), .C(_15665_), .Y(_15967_) );
	XOR2X1 XOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_15965_), .B(_15967_), .Y(_15968_) );
	XOR2X1 XOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_15968_), .B(_15960_), .Y(_15969_) );
	OAI21X1 OAI21X1_3384 ( .gnd(gnd), .vdd(vdd), .A(_15669_), .B(_15682_), .C(_15689_), .Y(_15970_) );
	INVX1 INVX1_2068 ( .gnd(gnd), .vdd(vdd), .A(_15970_), .Y(_15971_) );
	NOR2X1 NOR2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf3), .B(_14436_), .Y(_15972_) );
	NAND2X1 NAND2X1_3170 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf0), .B(aOperand_frameOut_24_bF_buf2), .Y(_15973_) );
	NAND2X1 NAND2X1_3171 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf0), .B(aOperand_frameOut_25_bF_buf3), .Y(_15974_) );
	XOR2X1 XOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_15973_), .B(_15974_), .Y(_15975_) );
	XOR2X1 XOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_15975_), .B(_15972_), .Y(_15976_) );
	NOR2X1 NOR2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_15349_), .B(_15673_), .Y(_15978_) );
	NOR2X1 NOR2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_15978_), .B(_15684_), .Y(_15979_) );
	NAND2X1 NAND2X1_3172 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf6), .B(aOperand_frameOut_28_), .Y(_15980_) );
	INVX1 INVX1_2069 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_28_), .Y(_15981_) );
	OAI21X1 OAI21X1_3385 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf1), .B(_15981_), .C(_15673_), .Y(_15982_) );
	OAI21X1 OAI21X1_3386 ( .gnd(gnd), .vdd(vdd), .A(_15675_), .B(_15980_), .C(_15982_), .Y(_15983_) );
	OAI21X1 OAI21X1_3387 ( .gnd(gnd), .vdd(vdd), .A(_12092_), .B(_15674_), .C(_15983_), .Y(_15984_) );
	NAND2X1 NAND2X1_3173 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf0), .B(aOperand_frameOut_26_), .Y(_15985_) );
	OR2X2 OR2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_15983_), .B(_15985_), .Y(_15986_) );
	NAND2X1 NAND2X1_3174 ( .gnd(gnd), .vdd(vdd), .A(_15984_), .B(_15986_), .Y(_15987_) );
	NAND2X1 NAND2X1_3175 ( .gnd(gnd), .vdd(vdd), .A(_15979_), .B(_15987_), .Y(_15989_) );
	OAI21X1 OAI21X1_3388 ( .gnd(gnd), .vdd(vdd), .A(_15349_), .B(_15673_), .C(_15680_), .Y(_15990_) );
	NAND3X1 NAND3X1_3363 ( .gnd(gnd), .vdd(vdd), .A(_15984_), .B(_15986_), .C(_15990_), .Y(_15991_) );
	AOI21X1 AOI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_15991_), .B(_15989_), .C(_15976_), .Y(_15992_) );
	INVX1 INVX1_2070 ( .gnd(gnd), .vdd(vdd), .A(_15976_), .Y(_15993_) );
	AND2X2 AND2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_15987_), .B(_15979_), .Y(_15994_) );
	NOR2X1 NOR2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_15979_), .B(_15987_), .Y(_15995_) );
	NOR3X1 NOR3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_15993_), .B(_15995_), .C(_15994_), .Y(_15996_) );
	OAI21X1 OAI21X1_3389 ( .gnd(gnd), .vdd(vdd), .A(_15992_), .B(_15996_), .C(_15971_), .Y(_15997_) );
	OAI21X1 OAI21X1_3390 ( .gnd(gnd), .vdd(vdd), .A(_15995_), .B(_15994_), .C(_15993_), .Y(_15998_) );
	NAND3X1 NAND3X1_3364 ( .gnd(gnd), .vdd(vdd), .A(_15976_), .B(_15989_), .C(_15991_), .Y(_16000_) );
	NAND3X1 NAND3X1_3365 ( .gnd(gnd), .vdd(vdd), .A(_15970_), .B(_16000_), .C(_15998_), .Y(_16001_) );
	AOI21X1 AOI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_15997_), .B(_16001_), .C(_15969_), .Y(_16002_) );
	XNOR2X1 XNOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_15968_), .B(_15960_), .Y(_16003_) );
	AOI21X1 AOI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_15998_), .B(_16000_), .C(_15970_), .Y(_16004_) );
	NOR3X1 NOR3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_15971_), .B(_15992_), .C(_15996_), .Y(_16005_) );
	NOR3X1 NOR3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_16004_), .B(_16003_), .C(_16005_), .Y(_16006_) );
	OAI21X1 OAI21X1_3391 ( .gnd(gnd), .vdd(vdd), .A(_16002_), .B(_16006_), .C(_15956_), .Y(_16007_) );
	OAI21X1 OAI21X1_3392 ( .gnd(gnd), .vdd(vdd), .A(_16004_), .B(_16005_), .C(_16003_), .Y(_16008_) );
	NAND3X1 NAND3X1_3366 ( .gnd(gnd), .vdd(vdd), .A(_15969_), .B(_16001_), .C(_15997_), .Y(_16009_) );
	NAND3X1 NAND3X1_3367 ( .gnd(gnd), .vdd(vdd), .A(_15954_), .B(_16009_), .C(_16008_), .Y(_16011_) );
	AOI21X1 AOI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_16007_), .B(_16011_), .C(_15953_), .Y(_16012_) );
	XOR2X1 XOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_15952_), .B(_15920_), .Y(_16013_) );
	AOI21X1 AOI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_16008_), .B(_16009_), .C(_15954_), .Y(_16014_) );
	NOR3X1 NOR3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_15956_), .B(_16002_), .C(_16006_), .Y(_16015_) );
	NOR3X1 NOR3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_16014_), .B(_16013_), .C(_16015_), .Y(_16016_) );
	OAI21X1 OAI21X1_3393 ( .gnd(gnd), .vdd(vdd), .A(_16012_), .B(_16016_), .C(_15919_), .Y(_16017_) );
	INVX1 INVX1_2071 ( .gnd(gnd), .vdd(vdd), .A(_15919_), .Y(_16018_) );
	OAI21X1 OAI21X1_3394 ( .gnd(gnd), .vdd(vdd), .A(_16014_), .B(_16015_), .C(_16013_), .Y(_16019_) );
	NAND3X1 NAND3X1_3368 ( .gnd(gnd), .vdd(vdd), .A(_16011_), .B(_15953_), .C(_16007_), .Y(_16020_) );
	NAND3X1 NAND3X1_3369 ( .gnd(gnd), .vdd(vdd), .A(_16020_), .B(_16019_), .C(_16018_), .Y(_16022_) );
	NAND3X1 NAND3X1_3370 ( .gnd(gnd), .vdd(vdd), .A(_16017_), .B(_16022_), .C(_15917_), .Y(_16023_) );
	NAND2X1 NAND2X1_3176 ( .gnd(gnd), .vdd(vdd), .A(_15912_), .B(_15916_), .Y(_16024_) );
	AOI21X1 AOI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_16019_), .B(_16020_), .C(_16018_), .Y(_16025_) );
	NOR3X1 NOR3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_15919_), .B(_16012_), .C(_16016_), .Y(_16026_) );
	OAI21X1 OAI21X1_3395 ( .gnd(gnd), .vdd(vdd), .A(_16025_), .B(_16026_), .C(_16024_), .Y(_16027_) );
	NAND3X1 NAND3X1_3371 ( .gnd(gnd), .vdd(vdd), .A(_15854_), .B(_16023_), .C(_16027_), .Y(_16028_) );
	AND2X2 AND2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_15723_), .B(_15717_), .Y(_16029_) );
	NOR3X1 NOR3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_16025_), .B(_16024_), .C(_16026_), .Y(_16030_) );
	AOI21X1 AOI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_16017_), .B(_16022_), .C(_15917_), .Y(_16031_) );
	OAI21X1 OAI21X1_3396 ( .gnd(gnd), .vdd(vdd), .A(_16031_), .B(_16030_), .C(_16029_), .Y(_16033_) );
	NAND3X1 NAND3X1_3372 ( .gnd(gnd), .vdd(vdd), .A(_16028_), .B(_16033_), .C(_15853_), .Y(_16034_) );
	NAND3X1 NAND3X1_3373 ( .gnd(gnd), .vdd(vdd), .A(_15794_), .B(_15843_), .C(_15848_), .Y(_16035_) );
	NAND3X1 NAND3X1_3374 ( .gnd(gnd), .vdd(vdd), .A(_15795_), .B(_15850_), .C(_15851_), .Y(_16036_) );
	NAND2X1 NAND2X1_3177 ( .gnd(gnd), .vdd(vdd), .A(_16035_), .B(_16036_), .Y(_16037_) );
	NOR3X1 NOR3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_16029_), .B(_16031_), .C(_16030_), .Y(_16038_) );
	AOI21X1 AOI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_16027_), .B(_16023_), .C(_15854_), .Y(_16039_) );
	OAI21X1 OAI21X1_3397 ( .gnd(gnd), .vdd(vdd), .A(_16039_), .B(_16038_), .C(_16037_), .Y(_16040_) );
	NAND3X1 NAND3X1_3375 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .B(_16034_), .C(_16040_), .Y(_16041_) );
	AND2X2 AND2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_15738_), .B(_15731_), .Y(_16042_) );
	OAI21X1 OAI21X1_3398 ( .gnd(gnd), .vdd(vdd), .A(_16031_), .B(_16030_), .C(_15854_), .Y(_16044_) );
	NAND3X1 NAND3X1_3376 ( .gnd(gnd), .vdd(vdd), .A(_16029_), .B(_16023_), .C(_16027_), .Y(_16045_) );
	AOI21X1 AOI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_16044_), .B(_16045_), .C(_16037_), .Y(_16046_) );
	AOI21X1 AOI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_16033_), .B(_16028_), .C(_15853_), .Y(_16047_) );
	OAI21X1 OAI21X1_3399 ( .gnd(gnd), .vdd(vdd), .A(_16046_), .B(_16047_), .C(_16042_), .Y(_16048_) );
	NAND3X1 NAND3X1_3377 ( .gnd(gnd), .vdd(vdd), .A(_15792_), .B(_16041_), .C(_16048_), .Y(_16049_) );
	INVX1 INVX1_2072 ( .gnd(gnd), .vdd(vdd), .A(_15792_), .Y(_16050_) );
	OAI21X1 OAI21X1_3400 ( .gnd(gnd), .vdd(vdd), .A(_16046_), .B(_16047_), .C(_15793_), .Y(_16051_) );
	NAND3X1 NAND3X1_3378 ( .gnd(gnd), .vdd(vdd), .A(_16042_), .B(_16034_), .C(_16040_), .Y(_16052_) );
	NAND3X1 NAND3X1_3379 ( .gnd(gnd), .vdd(vdd), .A(_16050_), .B(_16052_), .C(_16051_), .Y(_16053_) );
	NAND3X1 NAND3X1_3380 ( .gnd(gnd), .vdd(vdd), .A(_15791_), .B(_16049_), .C(_16053_), .Y(_16055_) );
	INVX1 INVX1_2073 ( .gnd(gnd), .vdd(vdd), .A(_15791_), .Y(_16056_) );
	AOI21X1 AOI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_16051_), .B(_16052_), .C(_16050_), .Y(_16057_) );
	AOI21X1 AOI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_16048_), .B(_16041_), .C(_15792_), .Y(_16058_) );
	OAI21X1 OAI21X1_3401 ( .gnd(gnd), .vdd(vdd), .A(_16057_), .B(_16058_), .C(_16056_), .Y(_16059_) );
	NAND3X1 NAND3X1_3381 ( .gnd(gnd), .vdd(vdd), .A(_15789_), .B(_16055_), .C(_16059_), .Y(_16060_) );
	OAI21X1 OAI21X1_3402 ( .gnd(gnd), .vdd(vdd), .A(_16057_), .B(_16058_), .C(_15791_), .Y(_16061_) );
	NAND3X1 NAND3X1_3382 ( .gnd(gnd), .vdd(vdd), .A(_16049_), .B(_16053_), .C(_16056_), .Y(_16062_) );
	NAND3X1 NAND3X1_3383 ( .gnd(gnd), .vdd(vdd), .A(_15757_), .B(_16062_), .C(_16061_), .Y(_16063_) );
	NAND2X1 NAND2X1_3178 ( .gnd(gnd), .vdd(vdd), .A(_16060_), .B(_16063_), .Y(_16064_) );
	XNOR2X1 XNOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .B(_16064_), .Y(mulOut_28_) );
	INVX1 INVX1_2074 ( .gnd(gnd), .vdd(vdd), .A(_16060_), .Y(_16066_) );
	AOI21X1 AOI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .B(_16063_), .C(_16066_), .Y(_16067_) );
	AOI21X1 AOI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_16040_), .B(_16034_), .C(_15793_), .Y(_16068_) );
	OAI21X1 OAI21X1_3403 ( .gnd(gnd), .vdd(vdd), .A(_16050_), .B(_16068_), .C(_16041_), .Y(_16069_) );
	NAND2X1 NAND2X1_3179 ( .gnd(gnd), .vdd(vdd), .A(_15843_), .B(_16035_), .Y(_16070_) );
	OAI21X1 OAI21X1_3404 ( .gnd(gnd), .vdd(vdd), .A(_16039_), .B(_16037_), .C(_16028_), .Y(_16071_) );
	NAND2X1 NAND2X1_3180 ( .gnd(gnd), .vdd(vdd), .A(_15832_), .B(_15838_), .Y(_16072_) );
	NOR2X1 NOR2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_15797_), .B(_15796_), .Y(_16073_) );
	NAND2X1 NAND2X1_3181 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf4), .B(adder_bOperand_29_), .Y(_16074_) );
	NAND2X1 NAND2X1_3182 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf0), .B(adder_bOperand_27_), .Y(_16076_) );
	XNOR2X1 XNOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_15797_), .B(_16076_), .Y(_16077_) );
	XOR2X1 XOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_16077_), .B(_16074_), .Y(_16078_) );
	OR2X2 OR2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_16078_), .B(_16073_), .Y(_16079_) );
	NAND2X1 NAND2X1_3183 ( .gnd(gnd), .vdd(vdd), .A(_16073_), .B(_16078_), .Y(_16080_) );
	NAND2X1 NAND2X1_3184 ( .gnd(gnd), .vdd(vdd), .A(_16080_), .B(_16079_), .Y(_16081_) );
	INVX1 INVX1_2075 ( .gnd(gnd), .vdd(vdd), .A(_16081_), .Y(_16082_) );
	INVX1 INVX1_2076 ( .gnd(gnd), .vdd(vdd), .A(_15827_), .Y(_16083_) );
	AOI21X1 AOI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_15804_), .B(_15829_), .C(_16083_), .Y(_16084_) );
	INVX1 INVX1_2077 ( .gnd(gnd), .vdd(vdd), .A(_16084_), .Y(_16085_) );
	NAND3X1 NAND3X1_3384 ( .gnd(gnd), .vdd(vdd), .A(_15805_), .B(_15819_), .C(_15816_), .Y(_16086_) );
	OAI21X1 OAI21X1_3405 ( .gnd(gnd), .vdd(vdd), .A(_15817_), .B(_15818_), .C(_16086_), .Y(_16087_) );
	OAI21X1 OAI21X1_3406 ( .gnd(gnd), .vdd(vdd), .A(_15807_), .B(_15808_), .C(_15814_), .Y(_16088_) );
	NAND2X1 NAND2X1_3185 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_5_bF_buf4), .B(adder_bOperand_24_), .Y(_16089_) );
	XNOR2X1 XNOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_15808_), .B(_16089_), .Y(_16090_) );
	OAI21X1 OAI21X1_3407 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_15806_), .C(_16090_), .Y(_16091_) );
	NAND2X1 NAND2X1_3186 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf1), .B(adder_bOperand_26_), .Y(_16092_) );
	OR2X2 OR2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_16090_), .B(_16092_), .Y(_16093_) );
	NAND2X1 NAND2X1_3187 ( .gnd(gnd), .vdd(vdd), .A(_16091_), .B(_16093_), .Y(_16094_) );
	NAND2X1 NAND2X1_3188 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf2), .B(adder_bOperand_22_bF_buf0), .Y(_16095_) );
	NAND2X1 NAND2X1_3189 ( .gnd(gnd), .vdd(vdd), .A(_15857_), .B(_15860_), .Y(_16098_) );
	OAI21X1 OAI21X1_3408 ( .gnd(gnd), .vdd(vdd), .A(_15519_), .B(_16095_), .C(_16098_), .Y(_16099_) );
	XNOR2X1 XNOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_16094_), .B(_16099_), .Y(_16100_) );
	XOR2X1 XOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_16100_), .B(_16088_), .Y(_16101_) );
	NAND3X1 NAND3X1_3385 ( .gnd(gnd), .vdd(vdd), .A(_15868_), .B(_15870_), .C(_15862_), .Y(_16102_) );
	NAND2X1 NAND2X1_3190 ( .gnd(gnd), .vdd(vdd), .A(_16102_), .B(_15873_), .Y(_16103_) );
	NAND2X1 NAND2X1_3191 ( .gnd(gnd), .vdd(vdd), .A(_16103_), .B(_16101_), .Y(_16104_) );
	XNOR2X1 XNOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_16100_), .B(_16088_), .Y(_16105_) );
	AND2X2 AND2X2_399 ( .gnd(gnd), .vdd(vdd), .A(_15873_), .B(_16102_), .Y(_16106_) );
	NAND2X1 NAND2X1_3192 ( .gnd(gnd), .vdd(vdd), .A(_16105_), .B(_16106_), .Y(_16107_) );
	NAND3X1 NAND3X1_3386 ( .gnd(gnd), .vdd(vdd), .A(_16087_), .B(_16104_), .C(_16107_), .Y(_16109_) );
	INVX1 INVX1_2078 ( .gnd(gnd), .vdd(vdd), .A(_16087_), .Y(_16110_) );
	NAND2X1 NAND2X1_3193 ( .gnd(gnd), .vdd(vdd), .A(_16101_), .B(_16106_), .Y(_16111_) );
	NAND2X1 NAND2X1_3194 ( .gnd(gnd), .vdd(vdd), .A(_16103_), .B(_16105_), .Y(_16112_) );
	NAND3X1 NAND3X1_3387 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_16112_), .C(_16111_), .Y(_16113_) );
	NAND3X1 NAND3X1_3388 ( .gnd(gnd), .vdd(vdd), .A(_16109_), .B(_16113_), .C(_16085_), .Y(_16114_) );
	AOI21X1 AOI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_16111_), .B(_16112_), .C(_16110_), .Y(_16115_) );
	INVX1 INVX1_2079 ( .gnd(gnd), .vdd(vdd), .A(_16113_), .Y(_16116_) );
	OAI21X1 OAI21X1_3409 ( .gnd(gnd), .vdd(vdd), .A(_16115_), .B(_16116_), .C(_16084_), .Y(_16117_) );
	NAND3X1 NAND3X1_3389 ( .gnd(gnd), .vdd(vdd), .A(_16082_), .B(_16114_), .C(_16117_), .Y(_16118_) );
	OAI21X1 OAI21X1_3410 ( .gnd(gnd), .vdd(vdd), .A(_16115_), .B(_16116_), .C(_16085_), .Y(_16120_) );
	NAND3X1 NAND3X1_3390 ( .gnd(gnd), .vdd(vdd), .A(_16109_), .B(_16084_), .C(_16113_), .Y(_16121_) );
	NAND3X1 NAND3X1_3391 ( .gnd(gnd), .vdd(vdd), .A(_16081_), .B(_16121_), .C(_16120_), .Y(_16122_) );
	NAND2X1 NAND2X1_3195 ( .gnd(gnd), .vdd(vdd), .A(_15906_), .B(_15912_), .Y(_16123_) );
	NAND3X1 NAND3X1_3392 ( .gnd(gnd), .vdd(vdd), .A(_16118_), .B(_16122_), .C(_16123_), .Y(_16124_) );
	AOI21X1 AOI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_16120_), .B(_16121_), .C(_16081_), .Y(_16125_) );
	AOI21X1 AOI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_16117_), .B(_16114_), .C(_16082_), .Y(_16126_) );
	INVX1 INVX1_2080 ( .gnd(gnd), .vdd(vdd), .A(_15906_), .Y(_16127_) );
	AOI21X1 AOI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_15855_), .B(_15910_), .C(_16127_), .Y(_16128_) );
	OAI21X1 OAI21X1_3411 ( .gnd(gnd), .vdd(vdd), .A(_16125_), .B(_16126_), .C(_16128_), .Y(_16129_) );
	NAND3X1 NAND3X1_3393 ( .gnd(gnd), .vdd(vdd), .A(_16072_), .B(_16124_), .C(_16129_), .Y(_16131_) );
	INVX1 INVX1_2081 ( .gnd(gnd), .vdd(vdd), .A(_16072_), .Y(_16132_) );
	NAND3X1 NAND3X1_3394 ( .gnd(gnd), .vdd(vdd), .A(_16128_), .B(_16118_), .C(_16122_), .Y(_16133_) );
	OAI21X1 OAI21X1_3412 ( .gnd(gnd), .vdd(vdd), .A(_16125_), .B(_16126_), .C(_16123_), .Y(_16134_) );
	NAND3X1 NAND3X1_3395 ( .gnd(gnd), .vdd(vdd), .A(_16133_), .B(_16132_), .C(_16134_), .Y(_16135_) );
	AND2X2 AND2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_16135_), .B(_16131_), .Y(_16136_) );
	AOI21X1 AOI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_15917_), .B(_16017_), .C(_16026_), .Y(_16137_) );
	OAI21X1 OAI21X1_3413 ( .gnd(gnd), .vdd(vdd), .A(_15895_), .B(_15897_), .C(_15899_), .Y(_16138_) );
	INVX1 INVX1_2082 ( .gnd(gnd), .vdd(vdd), .A(_16138_), .Y(_16139_) );
	NOR2X1 NOR2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_13294__bF_buf0), .B(_14564_), .Y(_16140_) );
	NAND2X1 NAND2X1_3196 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf2), .B(adder_bOperand_21_bF_buf3), .Y(_16142_) );
	XOR2X1 XOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_16095_), .B(_16142_), .Y(_16143_) );
	XOR2X1 XOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_16143_), .B(_16140_), .Y(_16144_) );
	OAI21X1 OAI21X1_3414 ( .gnd(gnd), .vdd(vdd), .A(_15531_), .B(_15863_), .C(_15870_), .Y(_16145_) );
	NAND2X1 NAND2X1_3197 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf2), .B(adder_bOperand_20_bF_buf2), .Y(_16146_) );
	NAND2X1 NAND2X1_3198 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf2), .B(adder_bOperand_19_bF_buf0), .Y(_16147_) );
	NAND2X1 NAND2X1_3199 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf1), .B(adder_bOperand_18_bF_buf0), .Y(_16148_) );
	OAI21X1 OAI21X1_3415 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_13067_), .C(_16148_), .Y(_16149_) );
	OAI21X1 OAI21X1_3416 ( .gnd(gnd), .vdd(vdd), .A(_15864_), .B(_16147_), .C(_16149_), .Y(_16150_) );
	XNOR2X1 XNOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_16150_), .B(_16146_), .Y(_16151_) );
	XNOR2X1 XNOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_16145_), .B(_16151_), .Y(_16153_) );
	XOR2X1 XOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_16153_), .B(_16144_), .Y(_16154_) );
	INVX1 INVX1_2083 ( .gnd(gnd), .vdd(vdd), .A(_16154_), .Y(_16155_) );
	OAI21X1 OAI21X1_3417 ( .gnd(gnd), .vdd(vdd), .A(_15896_), .B(_15892_), .C(_15890_), .Y(_16156_) );
	NAND2X1 NAND2X1_3200 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf0), .B(adder_bOperand_15_bF_buf2), .Y(_16157_) );
	OR2X2 OR2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_15550_), .B(_16157_), .Y(_16158_) );
	OAI21X1 OAI21X1_3418 ( .gnd(gnd), .vdd(vdd), .A(_15885_), .B(_15883_), .C(_16158_), .Y(_16159_) );
	INVX1 INVX1_2084 ( .gnd(gnd), .vdd(vdd), .A(_16159_), .Y(_16160_) );
	NAND2X1 NAND2X1_3201 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf2), .B(adder_bOperand_16_bF_buf1), .Y(_16161_) );
	NAND2X1 NAND2X1_3202 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf1), .B(adder_bOperand_15_bF_buf1), .Y(_16162_) );
	OAI21X1 OAI21X1_3419 ( .gnd(gnd), .vdd(vdd), .A(_11858_), .B(_12342_), .C(_16162_), .Y(_16164_) );
	OAI21X1 OAI21X1_3420 ( .gnd(gnd), .vdd(vdd), .A(_16157_), .B(_16161_), .C(_16164_), .Y(_16165_) );
	OAI21X1 OAI21X1_3421 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf3), .B(_12566_), .C(_16165_), .Y(_16166_) );
	NAND2X1 NAND2X1_3203 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf1), .B(adder_bOperand_17_bF_buf2), .Y(_16167_) );
	OR2X2 OR2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_16167_), .Y(_16168_) );
	NAND2X1 NAND2X1_3204 ( .gnd(gnd), .vdd(vdd), .A(_16166_), .B(_16168_), .Y(_16169_) );
	NAND2X1 NAND2X1_3205 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf3), .B(aOperand_frameOut_16_bF_buf1), .Y(_16170_) );
	NAND2X1 NAND2X1_3206 ( .gnd(gnd), .vdd(vdd), .A(_15921_), .B(_15925_), .Y(_16171_) );
	OAI21X1 OAI21X1_3422 ( .gnd(gnd), .vdd(vdd), .A(_15600_), .B(_16170_), .C(_16171_), .Y(_16172_) );
	XOR2X1 XOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_16169_), .B(_16172_), .Y(_16173_) );
	NOR2X1 NOR2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_16160_), .B(_16173_), .Y(_16175_) );
	XNOR2X1 XNOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_16169_), .B(_16172_), .Y(_16176_) );
	NOR2X1 NOR2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_16159_), .B(_16176_), .Y(_16177_) );
	OAI21X1 OAI21X1_3423 ( .gnd(gnd), .vdd(vdd), .A(_16177_), .B(_16175_), .C(_16156_), .Y(_16178_) );
	INVX1 INVX1_2085 ( .gnd(gnd), .vdd(vdd), .A(_15890_), .Y(_16179_) );
	AOI21X1 AOI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_15880_), .B(_15891_), .C(_16179_), .Y(_16180_) );
	NAND2X1 NAND2X1_3207 ( .gnd(gnd), .vdd(vdd), .A(_16159_), .B(_16176_), .Y(_16181_) );
	NAND2X1 NAND2X1_3208 ( .gnd(gnd), .vdd(vdd), .A(_16160_), .B(_16173_), .Y(_16182_) );
	NAND3X1 NAND3X1_3396 ( .gnd(gnd), .vdd(vdd), .A(_16181_), .B(_16180_), .C(_16182_), .Y(_16183_) );
	AOI21X1 AOI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_16178_), .B(_16183_), .C(_16155_), .Y(_16184_) );
	NAND3X1 NAND3X1_3397 ( .gnd(gnd), .vdd(vdd), .A(_16181_), .B(_16182_), .C(_16156_), .Y(_16186_) );
	OAI21X1 OAI21X1_3424 ( .gnd(gnd), .vdd(vdd), .A(_16177_), .B(_16175_), .C(_16180_), .Y(_16187_) );
	AOI21X1 AOI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_16187_), .B(_16186_), .C(_16154_), .Y(_16188_) );
	NAND3X1 NAND3X1_3398 ( .gnd(gnd), .vdd(vdd), .A(_15920_), .B(_15951_), .C(_15949_), .Y(_16189_) );
	AND2X2 AND2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_16189_), .B(_15951_), .Y(_16190_) );
	OAI21X1 OAI21X1_3425 ( .gnd(gnd), .vdd(vdd), .A(_16184_), .B(_16188_), .C(_16190_), .Y(_16191_) );
	NAND3X1 NAND3X1_3399 ( .gnd(gnd), .vdd(vdd), .A(_16154_), .B(_16186_), .C(_16187_), .Y(_16192_) );
	NAND3X1 NAND3X1_3400 ( .gnd(gnd), .vdd(vdd), .A(_16183_), .B(_16178_), .C(_16155_), .Y(_16193_) );
	NAND2X1 NAND2X1_3209 ( .gnd(gnd), .vdd(vdd), .A(_15951_), .B(_16189_), .Y(_16194_) );
	NAND3X1 NAND3X1_3401 ( .gnd(gnd), .vdd(vdd), .A(_16192_), .B(_16194_), .C(_16193_), .Y(_16195_) );
	NAND2X1 NAND2X1_3210 ( .gnd(gnd), .vdd(vdd), .A(_16195_), .B(_16191_), .Y(_16197_) );
	NAND2X1 NAND2X1_3211 ( .gnd(gnd), .vdd(vdd), .A(_16139_), .B(_16197_), .Y(_16198_) );
	NAND3X1 NAND3X1_3402 ( .gnd(gnd), .vdd(vdd), .A(_16195_), .B(_16138_), .C(_16191_), .Y(_16199_) );
	AND2X2 AND2X2_402 ( .gnd(gnd), .vdd(vdd), .A(_16198_), .B(_16199_), .Y(_16200_) );
	AOI21X1 AOI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_16007_), .B(_15953_), .C(_16015_), .Y(_16201_) );
	OAI21X1 OAI21X1_3426 ( .gnd(gnd), .vdd(vdd), .A(_15937_), .B(_15940_), .C(_15942_), .Y(_16202_) );
	NAND2X1 NAND2X1_3212 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf0), .B(aOperand_frameOut_15_bF_buf2), .Y(_16203_) );
	NAND2X1 NAND2X1_3213 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf2), .B(aOperand_frameOut_17_bF_buf0), .Y(_16204_) );
	XOR2X1 XOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_16170_), .B(_16204_), .Y(_16205_) );
	XNOR2X1 XNOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_16205_), .B(_16203_), .Y(_16206_) );
	OAI21X1 OAI21X1_3427 ( .gnd(gnd), .vdd(vdd), .A(_15927_), .B(_15931_), .C(_15939_), .Y(_16208_) );
	NAND2X1 NAND2X1_3214 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf4), .B(aOperand_frameOut_19_bF_buf0), .Y(_16209_) );
	NAND2X1 NAND2X1_3215 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf1), .B(aOperand_frameOut_20_bF_buf2), .Y(_16210_) );
	NAND2X1 NAND2X1_3216 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf3), .B(aOperand_frameOut_20_bF_buf1), .Y(_16211_) );
	OAI21X1 OAI21X1_3428 ( .gnd(gnd), .vdd(vdd), .A(_16887_), .B(_13224_), .C(_16211_), .Y(_16212_) );
	OAI21X1 OAI21X1_3429 ( .gnd(gnd), .vdd(vdd), .A(_16209_), .B(_16210_), .C(_16212_), .Y(_16213_) );
	OAI21X1 OAI21X1_3430 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf3), .B(_13796_), .C(_16213_), .Y(_16214_) );
	NAND2X1 NAND2X1_3217 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf3), .B(aOperand_frameOut_18_bF_buf3), .Y(_16215_) );
	OR2X2 OR2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_16215_), .Y(_16216_) );
	NAND2X1 NAND2X1_3218 ( .gnd(gnd), .vdd(vdd), .A(_16214_), .B(_16216_), .Y(_16217_) );
	XNOR2X1 XNOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_16208_), .B(_16217_), .Y(_16219_) );
	NAND2X1 NAND2X1_3219 ( .gnd(gnd), .vdd(vdd), .A(_16206_), .B(_16219_), .Y(_16220_) );
	INVX1 INVX1_2086 ( .gnd(gnd), .vdd(vdd), .A(_16206_), .Y(_16221_) );
	XOR2X1 XOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_16208_), .B(_16217_), .Y(_16222_) );
	NAND2X1 NAND2X1_3220 ( .gnd(gnd), .vdd(vdd), .A(_16221_), .B(_16222_), .Y(_16223_) );
	NOR2X1 NOR2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_15967_), .B(_15965_), .Y(_16224_) );
	AOI21X1 AOI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_15968_), .B(_15960_), .C(_16224_), .Y(_16225_) );
	INVX1 INVX1_2087 ( .gnd(gnd), .vdd(vdd), .A(_16225_), .Y(_16226_) );
	NAND3X1 NAND3X1_3403 ( .gnd(gnd), .vdd(vdd), .A(_16220_), .B(_16223_), .C(_16226_), .Y(_16227_) );
	NOR2X1 NOR2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_16221_), .B(_16222_), .Y(_16228_) );
	NOR2X1 NOR2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_16206_), .B(_16219_), .Y(_16230_) );
	OAI21X1 OAI21X1_3431 ( .gnd(gnd), .vdd(vdd), .A(_16230_), .B(_16228_), .C(_16225_), .Y(_16231_) );
	NAND3X1 NAND3X1_3404 ( .gnd(gnd), .vdd(vdd), .A(_16202_), .B(_16231_), .C(_16227_), .Y(_16232_) );
	INVX1 INVX1_2088 ( .gnd(gnd), .vdd(vdd), .A(_16202_), .Y(_16233_) );
	NAND3X1 NAND3X1_3405 ( .gnd(gnd), .vdd(vdd), .A(_16225_), .B(_16220_), .C(_16223_), .Y(_16234_) );
	OAI21X1 OAI21X1_3432 ( .gnd(gnd), .vdd(vdd), .A(_16230_), .B(_16228_), .C(_16226_), .Y(_16235_) );
	NAND3X1 NAND3X1_3406 ( .gnd(gnd), .vdd(vdd), .A(_16233_), .B(_16234_), .C(_16235_), .Y(_16236_) );
	AND2X2 AND2X2_403 ( .gnd(gnd), .vdd(vdd), .A(_16232_), .B(_16236_), .Y(_16237_) );
	AOI21X1 AOI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_15997_), .B(_15969_), .C(_16005_), .Y(_16238_) );
	NAND2X1 NAND2X1_3221 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf1), .B(aOperand_frameOut_22_bF_buf0), .Y(_16239_) );
	NOR2X1 NOR2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_15648_), .B(_16239_), .Y(_16241_) );
	NOR2X1 NOR2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_15961_), .B(_15964_), .Y(_16242_) );
	NOR2X1 NOR2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_16241_), .B(_16242_), .Y(_16243_) );
	INVX1 INVX1_2089 ( .gnd(gnd), .vdd(vdd), .A(_16243_), .Y(_16244_) );
	NAND2X1 NAND2X1_3222 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf0), .B(aOperand_frameOut_23_), .Y(_16245_) );
	NAND2X1 NAND2X1_3223 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf0), .B(aOperand_frameOut_23_), .Y(_16246_) );
	OAI21X1 OAI21X1_3433 ( .gnd(gnd), .vdd(vdd), .A(_13830_), .B(_14125_), .C(_16246_), .Y(_16247_) );
	OAI21X1 OAI21X1_3434 ( .gnd(gnd), .vdd(vdd), .A(_16239_), .B(_16245_), .C(_16247_), .Y(_16248_) );
	OAI21X1 OAI21X1_3435 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf3), .B(_13812_), .C(_16248_), .Y(_16249_) );
	NAND2X1 NAND2X1_3224 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf3), .B(aOperand_frameOut_21_bF_buf1), .Y(_16250_) );
	OR2X2 OR2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_16248_), .B(_16250_), .Y(_16252_) );
	NAND2X1 NAND2X1_3225 ( .gnd(gnd), .vdd(vdd), .A(_16249_), .B(_16252_), .Y(_16253_) );
	NAND2X1 NAND2X1_3226 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf5), .B(aOperand_frameOut_25_bF_buf2), .Y(_16254_) );
	NAND2X1 NAND2X1_3227 ( .gnd(gnd), .vdd(vdd), .A(_15972_), .B(_15975_), .Y(_16255_) );
	OAI21X1 OAI21X1_3436 ( .gnd(gnd), .vdd(vdd), .A(_15663_), .B(_16254_), .C(_16255_), .Y(_16256_) );
	NOR2X1 NOR2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_16256_), .B(_16253_), .Y(_16257_) );
	AND2X2 AND2X2_404 ( .gnd(gnd), .vdd(vdd), .A(_16253_), .B(_16256_), .Y(_16258_) );
	OAI21X1 OAI21X1_3437 ( .gnd(gnd), .vdd(vdd), .A(_16257_), .B(_16258_), .C(_16244_), .Y(_16259_) );
	NOR2X1 NOR2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_16257_), .B(_16258_), .Y(_16260_) );
	NAND2X1 NAND2X1_3228 ( .gnd(gnd), .vdd(vdd), .A(_16243_), .B(_16260_), .Y(_16261_) );
	AND2X2 AND2X2_405 ( .gnd(gnd), .vdd(vdd), .A(_16261_), .B(_16259_), .Y(_16263_) );
	AOI21X1 AOI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_15976_), .B(_15989_), .C(_15995_), .Y(_16264_) );
	NAND2X1 NAND2X1_3229 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf3), .B(aOperand_frameOut_24_bF_buf1), .Y(_16265_) );
	NAND2X1 NAND2X1_3230 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf5), .B(aOperand_frameOut_26_), .Y(_16266_) );
	XOR2X1 XOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_16254_), .B(_16266_), .Y(_16267_) );
	XNOR2X1 XNOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_16267_), .B(_16265_), .Y(_16268_) );
	NAND2X1 NAND2X1_3231 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf3), .B(aOperand_frameOut_28_), .Y(_16269_) );
	NOR2X1 NOR2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_15673_), .B(_16269_), .Y(_16270_) );
	NOR2X1 NOR2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_15985_), .B(_15983_), .Y(_16271_) );
	NOR2X1 NOR2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_16270_), .B(_16271_), .Y(_16272_) );
	NAND2X1 NAND2X1_3232 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf5), .B(aOperand_frameOut_27_), .Y(_16274_) );
	NAND2X1 NAND2X1_3233 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf5), .B(aOperand_frameOut_29_), .Y(_16275_) );
	NAND2X1 NAND2X1_3234 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf2), .B(aOperand_frameOut_29_), .Y(_16276_) );
	OAI21X1 OAI21X1_3438 ( .gnd(gnd), .vdd(vdd), .A(_11776__bF_buf1), .B(_15981_), .C(_16276_), .Y(_16277_) );
	OAI21X1 OAI21X1_3439 ( .gnd(gnd), .vdd(vdd), .A(_16269_), .B(_16275_), .C(_16277_), .Y(_16278_) );
	XNOR2X1 XNOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_16278_), .B(_16274_), .Y(_16279_) );
	NAND2X1 NAND2X1_3235 ( .gnd(gnd), .vdd(vdd), .A(_16279_), .B(_16272_), .Y(_16280_) );
	XOR2X1 XOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_16278_), .B(_16274_), .Y(_16281_) );
	OAI21X1 OAI21X1_3440 ( .gnd(gnd), .vdd(vdd), .A(_16270_), .B(_16271_), .C(_16281_), .Y(_16282_) );
	AOI21X1 AOI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_16280_), .B(_16282_), .C(_16268_), .Y(_16283_) );
	INVX1 INVX1_2090 ( .gnd(gnd), .vdd(vdd), .A(_16268_), .Y(_16285_) );
	NAND2X1 NAND2X1_3236 ( .gnd(gnd), .vdd(vdd), .A(_16282_), .B(_16280_), .Y(_16286_) );
	NOR2X1 NOR2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_16285_), .B(_16286_), .Y(_16287_) );
	OAI21X1 OAI21X1_3441 ( .gnd(gnd), .vdd(vdd), .A(_16283_), .B(_16287_), .C(_16264_), .Y(_16288_) );
	INVX1 INVX1_2091 ( .gnd(gnd), .vdd(vdd), .A(_16264_), .Y(_16289_) );
	INVX1 INVX1_2092 ( .gnd(gnd), .vdd(vdd), .A(_16283_), .Y(_16290_) );
	OR2X2 OR2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_16286_), .B(_16285_), .Y(_16291_) );
	NAND3X1 NAND3X1_3407 ( .gnd(gnd), .vdd(vdd), .A(_16290_), .B(_16289_), .C(_16291_), .Y(_16292_) );
	AOI21X1 AOI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_16292_), .B(_16288_), .C(_16263_), .Y(_16293_) );
	NAND2X1 NAND2X1_3237 ( .gnd(gnd), .vdd(vdd), .A(_16259_), .B(_16261_), .Y(_16294_) );
	AOI21X1 AOI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_16291_), .B(_16290_), .C(_16289_), .Y(_16296_) );
	NOR3X1 NOR3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_16264_), .B(_16283_), .C(_16287_), .Y(_16297_) );
	NOR3X1 NOR3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_16294_), .B(_16297_), .C(_16296_), .Y(_16298_) );
	OAI21X1 OAI21X1_3442 ( .gnd(gnd), .vdd(vdd), .A(_16293_), .B(_16298_), .C(_16238_), .Y(_16299_) );
	INVX1 INVX1_2093 ( .gnd(gnd), .vdd(vdd), .A(_16238_), .Y(_16300_) );
	OAI21X1 OAI21X1_3443 ( .gnd(gnd), .vdd(vdd), .A(_16297_), .B(_16296_), .C(_16294_), .Y(_16301_) );
	NAND3X1 NAND3X1_3408 ( .gnd(gnd), .vdd(vdd), .A(_16288_), .B(_16292_), .C(_16263_), .Y(_16302_) );
	NAND3X1 NAND3X1_3409 ( .gnd(gnd), .vdd(vdd), .A(_16301_), .B(_16302_), .C(_16300_), .Y(_16303_) );
	AOI21X1 AOI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_16299_), .B(_16303_), .C(_16237_), .Y(_16304_) );
	NAND2X1 NAND2X1_3238 ( .gnd(gnd), .vdd(vdd), .A(_16236_), .B(_16232_), .Y(_16305_) );
	AOI21X1 AOI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_16301_), .B(_16302_), .C(_16300_), .Y(_16307_) );
	NOR3X1 NOR3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_16238_), .B(_16293_), .C(_16298_), .Y(_16308_) );
	NOR3X1 NOR3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_16305_), .B(_16307_), .C(_16308_), .Y(_16309_) );
	OAI21X1 OAI21X1_3444 ( .gnd(gnd), .vdd(vdd), .A(_16304_), .B(_16309_), .C(_16201_), .Y(_16310_) );
	OAI21X1 OAI21X1_3445 ( .gnd(gnd), .vdd(vdd), .A(_16014_), .B(_16013_), .C(_16011_), .Y(_16311_) );
	OAI21X1 OAI21X1_3446 ( .gnd(gnd), .vdd(vdd), .A(_16307_), .B(_16308_), .C(_16305_), .Y(_16312_) );
	NAND3X1 NAND3X1_3410 ( .gnd(gnd), .vdd(vdd), .A(_16303_), .B(_16299_), .C(_16237_), .Y(_16313_) );
	NAND3X1 NAND3X1_3411 ( .gnd(gnd), .vdd(vdd), .A(_16311_), .B(_16313_), .C(_16312_), .Y(_16314_) );
	AOI21X1 AOI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_16310_), .B(_16314_), .C(_16200_), .Y(_16315_) );
	NAND2X1 NAND2X1_3239 ( .gnd(gnd), .vdd(vdd), .A(_16199_), .B(_16198_), .Y(_16316_) );
	AOI21X1 AOI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_16312_), .B(_16313_), .C(_16311_), .Y(_16318_) );
	NOR3X1 NOR3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_16201_), .B(_16304_), .C(_16309_), .Y(_16319_) );
	NOR3X1 NOR3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_16318_), .B(_16316_), .C(_16319_), .Y(_16320_) );
	OAI21X1 OAI21X1_3447 ( .gnd(gnd), .vdd(vdd), .A(_16315_), .B(_16320_), .C(_16137_), .Y(_16321_) );
	OAI21X1 OAI21X1_3448 ( .gnd(gnd), .vdd(vdd), .A(_16025_), .B(_16024_), .C(_16022_), .Y(_16322_) );
	OAI21X1 OAI21X1_3449 ( .gnd(gnd), .vdd(vdd), .A(_16318_), .B(_16319_), .C(_16316_), .Y(_16323_) );
	NAND3X1 NAND3X1_3412 ( .gnd(gnd), .vdd(vdd), .A(_16314_), .B(_16310_), .C(_16200_), .Y(_16324_) );
	NAND3X1 NAND3X1_3413 ( .gnd(gnd), .vdd(vdd), .A(_16322_), .B(_16324_), .C(_16323_), .Y(_16325_) );
	NAND3X1 NAND3X1_3414 ( .gnd(gnd), .vdd(vdd), .A(_16321_), .B(_16325_), .C(_16136_), .Y(_16326_) );
	NAND2X1 NAND2X1_3240 ( .gnd(gnd), .vdd(vdd), .A(_16131_), .B(_16135_), .Y(_16327_) );
	AOI21X1 AOI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_16323_), .B(_16324_), .C(_16322_), .Y(_16329_) );
	NOR3X1 NOR3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_16137_), .B(_16315_), .C(_16320_), .Y(_16330_) );
	OAI21X1 OAI21X1_3450 ( .gnd(gnd), .vdd(vdd), .A(_16329_), .B(_16330_), .C(_16327_), .Y(_16331_) );
	NAND3X1 NAND3X1_3415 ( .gnd(gnd), .vdd(vdd), .A(_16071_), .B(_16331_), .C(_16326_), .Y(_16332_) );
	AOI21X1 AOI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_15853_), .B(_16033_), .C(_16038_), .Y(_16333_) );
	OAI21X1 OAI21X1_3451 ( .gnd(gnd), .vdd(vdd), .A(_16329_), .B(_16330_), .C(_16136_), .Y(_16334_) );
	NAND3X1 NAND3X1_3416 ( .gnd(gnd), .vdd(vdd), .A(_16325_), .B(_16321_), .C(_16327_), .Y(_16335_) );
	NAND3X1 NAND3X1_3417 ( .gnd(gnd), .vdd(vdd), .A(_16333_), .B(_16335_), .C(_16334_), .Y(_16336_) );
	NAND3X1 NAND3X1_3418 ( .gnd(gnd), .vdd(vdd), .A(_16070_), .B(_16336_), .C(_16332_), .Y(_16337_) );
	INVX1 INVX1_2094 ( .gnd(gnd), .vdd(vdd), .A(_16070_), .Y(_16338_) );
	AOI21X1 AOI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_16334_), .B(_16335_), .C(_16333_), .Y(_16340_) );
	AOI21X1 AOI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_16326_), .B(_16331_), .C(_16071_), .Y(_16341_) );
	OAI21X1 OAI21X1_3452 ( .gnd(gnd), .vdd(vdd), .A(_16340_), .B(_16341_), .C(_16338_), .Y(_16342_) );
	NAND3X1 NAND3X1_3419 ( .gnd(gnd), .vdd(vdd), .A(_16069_), .B(_16337_), .C(_16342_), .Y(_16343_) );
	NOR3X1 NOR3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_16042_), .B(_16046_), .C(_16047_), .Y(_16344_) );
	AOI21X1 AOI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_15792_), .B(_16048_), .C(_16344_), .Y(_16345_) );
	OAI21X1 OAI21X1_3453 ( .gnd(gnd), .vdd(vdd), .A(_16340_), .B(_16341_), .C(_16070_), .Y(_16346_) );
	NAND3X1 NAND3X1_3420 ( .gnd(gnd), .vdd(vdd), .A(_16338_), .B(_16336_), .C(_16332_), .Y(_16347_) );
	NAND3X1 NAND3X1_3421 ( .gnd(gnd), .vdd(vdd), .A(_16345_), .B(_16347_), .C(_16346_), .Y(_16348_) );
	NAND3X1 NAND3X1_3422 ( .gnd(gnd), .vdd(vdd), .A(_16055_), .B(_16343_), .C(_16348_), .Y(_16349_) );
	INVX1 INVX1_2095 ( .gnd(gnd), .vdd(vdd), .A(_16055_), .Y(_16351_) );
	NAND3X1 NAND3X1_3423 ( .gnd(gnd), .vdd(vdd), .A(_16345_), .B(_16337_), .C(_16342_), .Y(_16352_) );
	NAND3X1 NAND3X1_3424 ( .gnd(gnd), .vdd(vdd), .A(_16069_), .B(_16347_), .C(_16346_), .Y(_16353_) );
	NAND3X1 NAND3X1_3425 ( .gnd(gnd), .vdd(vdd), .A(_16352_), .B(_16353_), .C(_16351_), .Y(_16354_) );
	NAND2X1 NAND2X1_3241 ( .gnd(gnd), .vdd(vdd), .A(_16349_), .B(_16354_), .Y(_16355_) );
	XNOR2X1 XNOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_16067_), .B(_16355_), .Y(mulOut_29_) );
	AND2X2 AND2X2_406 ( .gnd(gnd), .vdd(vdd), .A(_14530_), .B(_13925_), .Y(_16356_) );
	NAND2X1 NAND2X1_3242 ( .gnd(gnd), .vdd(vdd), .A(_16356_), .B(_13916_), .Y(_16357_) );
	AOI21X1 AOI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_14221_), .B(_14220_), .C(_13899_), .Y(_16358_) );
	AOI21X1 AOI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_14215_), .B(_14218_), .C(_13893_), .Y(_16359_) );
	NAND2X1 NAND2X1_3243 ( .gnd(gnd), .vdd(vdd), .A(_14216_), .B(_14217_), .Y(_16361_) );
	AOI22X1 AOI22X1_372 ( .gnd(gnd), .vdd(vdd), .A(_13930_), .B(_16361_), .C(_14526_), .D(_14527_), .Y(_16362_) );
	AOI21X1 AOI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_14523_), .B(_14517_), .C(_14215_), .Y(_16363_) );
	OAI22X1 OAI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(_16358_), .B(_16359_), .C(_16362_), .D(_16363_), .Y(_16364_) );
	NAND2X1 NAND2X1_3244 ( .gnd(gnd), .vdd(vdd), .A(_14534_), .B(_14536_), .Y(_16365_) );
	OAI21X1 OAI21X1_3454 ( .gnd(gnd), .vdd(vdd), .A(_13907_), .B(_16364_), .C(_16365_), .Y(_16366_) );
	AOI21X1 AOI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_13924_), .B(_16356_), .C(_16366_), .Y(_16367_) );
	AOI21X1 AOI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_16367_), .B(_16357_), .C(_15778_), .Y(_16368_) );
	INVX1 INVX1_2096 ( .gnd(gnd), .vdd(vdd), .A(_15773_), .Y(_16369_) );
	AOI21X1 AOI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_15442_), .B(_15774_), .C(_16369_), .Y(_16370_) );
	OAI21X1 OAI21X1_3455 ( .gnd(gnd), .vdd(vdd), .A(_15784_), .B(_15125_), .C(_16370_), .Y(_16372_) );
	AOI21X1 AOI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_16349_), .B(_16354_), .C(_16064_), .Y(_16373_) );
	OAI21X1 OAI21X1_3456 ( .gnd(gnd), .vdd(vdd), .A(_16372_), .B(_16368_), .C(_16373_), .Y(_16374_) );
	AOI21X1 AOI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_16352_), .B(_16353_), .C(_16055_), .Y(_16375_) );
	AOI21X1 AOI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_16355_), .B(_16066_), .C(_16375_), .Y(_16376_) );
	OAI21X1 OAI21X1_3457 ( .gnd(gnd), .vdd(vdd), .A(_16338_), .B(_16341_), .C(_16332_), .Y(_16377_) );
	NAND2X1 NAND2X1_3245 ( .gnd(gnd), .vdd(vdd), .A(_16124_), .B(_16131_), .Y(_16378_) );
	OAI21X1 OAI21X1_3458 ( .gnd(gnd), .vdd(vdd), .A(_16329_), .B(_16327_), .C(_16325_), .Y(_16379_) );
	INVX1 INVX1_2097 ( .gnd(gnd), .vdd(vdd), .A(_16379_), .Y(_16380_) );
	NAND2X1 NAND2X1_3246 ( .gnd(gnd), .vdd(vdd), .A(_16114_), .B(_16118_), .Y(_16381_) );
	NAND2X1 NAND2X1_3247 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf3), .B(adder_bOperand_30_), .Y(_16383_) );
	NOR2X1 NOR2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_15797_), .B(_16076_), .Y(_16384_) );
	NOR2X1 NOR2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_16074_), .B(_16077_), .Y(_16385_) );
	NOR2X1 NOR2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_16384_), .B(_16385_), .Y(_16386_) );
	NAND2X1 NAND2X1_3248 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf1), .B(adder_bOperand_29_), .Y(_16387_) );
	NAND2X1 NAND2X1_3249 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_3_bF_buf0), .B(adder_bOperand_28_), .Y(_16388_) );
	OAI22X1 OAI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_12310__bF_buf0), .B(_15798_), .C(_12048_), .D(_15454_), .Y(_16389_) );
	OAI21X1 OAI21X1_3459 ( .gnd(gnd), .vdd(vdd), .A(_16076_), .B(_16388_), .C(_16389_), .Y(_16390_) );
	NAND2X1 NAND2X1_3250 ( .gnd(gnd), .vdd(vdd), .A(_16387_), .B(_16390_), .Y(_16391_) );
	OR2X2 OR2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_16390_), .B(_16387_), .Y(_16392_) );
	NAND2X1 NAND2X1_3251 ( .gnd(gnd), .vdd(vdd), .A(_16391_), .B(_16392_), .Y(_16393_) );
	OR2X2 OR2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_16386_), .B(_16393_), .Y(_16394_) );
	NAND2X1 NAND2X1_3252 ( .gnd(gnd), .vdd(vdd), .A(_16393_), .B(_16386_), .Y(_16395_) );
	NAND2X1 NAND2X1_3253 ( .gnd(gnd), .vdd(vdd), .A(_16395_), .B(_16394_), .Y(_16396_) );
	XNOR2X1 XNOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_16396_), .B(_16383_), .Y(_16397_) );
	NAND2X1 NAND2X1_3254 ( .gnd(gnd), .vdd(vdd), .A(_16080_), .B(_16397_), .Y(_16398_) );
	NOR2X1 NOR2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_16080_), .B(_16397_), .Y(_16399_) );
	INVX1 INVX1_2098 ( .gnd(gnd), .vdd(vdd), .A(_16399_), .Y(_16400_) );
	NAND2X1 NAND2X1_3255 ( .gnd(gnd), .vdd(vdd), .A(_16398_), .B(_16400_), .Y(_16401_) );
	OAI21X1 OAI21X1_3460 ( .gnd(gnd), .vdd(vdd), .A(_16105_), .B(_16106_), .C(_16109_), .Y(_16402_) );
	NAND3X1 NAND3X1_3426 ( .gnd(gnd), .vdd(vdd), .A(_16091_), .B(_16093_), .C(_16099_), .Y(_16404_) );
	NAND2X1 NAND2X1_3256 ( .gnd(gnd), .vdd(vdd), .A(_16088_), .B(_16100_), .Y(_16405_) );
	NAND2X1 NAND2X1_3257 ( .gnd(gnd), .vdd(vdd), .A(_16404_), .B(_16405_), .Y(_16406_) );
	INVX1 INVX1_2099 ( .gnd(gnd), .vdd(vdd), .A(_16406_), .Y(_16407_) );
	OAI21X1 OAI21X1_3461 ( .gnd(gnd), .vdd(vdd), .A(_15808_), .B(_16089_), .C(_16093_), .Y(_16408_) );
	NAND2X1 NAND2X1_3258 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf4), .B(adder_bOperand_26_), .Y(_16409_) );
	NAND2X1 NAND2X1_3259 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_6_bF_buf0), .B(adder_bOperand_25_), .Y(_16410_) );
	OAI22X1 OAI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_14827_), .C(_13294__bF_buf3), .D(_14544_), .Y(_16411_) );
	OAI21X1 OAI21X1_3462 ( .gnd(gnd), .vdd(vdd), .A(_16089_), .B(_16410_), .C(_16411_), .Y(_16412_) );
	XNOR2X1 XNOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_16412_), .B(_16409_), .Y(_16413_) );
	NAND2X1 NAND2X1_3260 ( .gnd(gnd), .vdd(vdd), .A(_16140_), .B(_16143_), .Y(_16416_) );
	OAI21X1 OAI21X1_3463 ( .gnd(gnd), .vdd(vdd), .A(_16095_), .B(_16142_), .C(_16416_), .Y(_16417_) );
	XNOR2X1 XNOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_16417_), .B(_16413_), .Y(_16418_) );
	XNOR2X1 XNOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_16418_), .B(_16408_), .Y(_16419_) );
	OAI21X1 OAI21X1_3464 ( .gnd(gnd), .vdd(vdd), .A(_15812__bF_buf3), .B(_13334_), .C(_16150_), .Y(_16420_) );
	OR2X2 OR2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_16150_), .B(_16146_), .Y(_16421_) );
	NAND3X1 NAND3X1_3427 ( .gnd(gnd), .vdd(vdd), .A(_16420_), .B(_16421_), .C(_16145_), .Y(_16422_) );
	NAND2X1 NAND2X1_3261 ( .gnd(gnd), .vdd(vdd), .A(_16144_), .B(_16153_), .Y(_16423_) );
	NAND2X1 NAND2X1_3262 ( .gnd(gnd), .vdd(vdd), .A(_16422_), .B(_16423_), .Y(_16424_) );
	XOR2X1 XOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_16419_), .B(_16424_), .Y(_16425_) );
	NAND2X1 NAND2X1_3263 ( .gnd(gnd), .vdd(vdd), .A(_16407_), .B(_16425_), .Y(_16427_) );
	NAND3X1 NAND3X1_3428 ( .gnd(gnd), .vdd(vdd), .A(_16422_), .B(_16423_), .C(_16419_), .Y(_16428_) );
	AND2X2 AND2X2_407 ( .gnd(gnd), .vdd(vdd), .A(_16423_), .B(_16422_), .Y(_16429_) );
	OR2X2 OR2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_16429_), .B(_16419_), .Y(_16430_) );
	NAND3X1 NAND3X1_3429 ( .gnd(gnd), .vdd(vdd), .A(_16406_), .B(_16428_), .C(_16430_), .Y(_16431_) );
	NAND2X1 NAND2X1_3264 ( .gnd(gnd), .vdd(vdd), .A(_16431_), .B(_16427_), .Y(_16432_) );
	XOR2X1 XOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_16432_), .B(_16402_), .Y(_16433_) );
	OR2X2 OR2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_16433_), .B(_16401_), .Y(_16434_) );
	NAND2X1 NAND2X1_3265 ( .gnd(gnd), .vdd(vdd), .A(_16401_), .B(_16433_), .Y(_16435_) );
	OAI21X1 OAI21X1_3465 ( .gnd(gnd), .vdd(vdd), .A(_16139_), .B(_16197_), .C(_16195_), .Y(_16436_) );
	NAND3X1 NAND3X1_3430 ( .gnd(gnd), .vdd(vdd), .A(_16435_), .B(_16436_), .C(_16434_), .Y(_16438_) );
	NOR2X1 NOR2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_16401_), .B(_16433_), .Y(_16439_) );
	AND2X2 AND2X2_408 ( .gnd(gnd), .vdd(vdd), .A(_16433_), .B(_16401_), .Y(_16440_) );
	INVX1 INVX1_2100 ( .gnd(gnd), .vdd(vdd), .A(_16436_), .Y(_16441_) );
	OAI21X1 OAI21X1_3466 ( .gnd(gnd), .vdd(vdd), .A(_16439_), .B(_16440_), .C(_16441_), .Y(_16442_) );
	NAND3X1 NAND3X1_3431 ( .gnd(gnd), .vdd(vdd), .A(_16381_), .B(_16438_), .C(_16442_), .Y(_16443_) );
	INVX1 INVX1_2101 ( .gnd(gnd), .vdd(vdd), .A(_16381_), .Y(_16444_) );
	OAI21X1 OAI21X1_3467 ( .gnd(gnd), .vdd(vdd), .A(_16439_), .B(_16440_), .C(_16436_), .Y(_16445_) );
	NAND3X1 NAND3X1_3432 ( .gnd(gnd), .vdd(vdd), .A(_16435_), .B(_16441_), .C(_16434_), .Y(_16446_) );
	NAND3X1 NAND3X1_3433 ( .gnd(gnd), .vdd(vdd), .A(_16444_), .B(_16446_), .C(_16445_), .Y(_16447_) );
	NAND2X1 NAND2X1_3266 ( .gnd(gnd), .vdd(vdd), .A(_16443_), .B(_16447_), .Y(_16449_) );
	NAND2X1 NAND2X1_3267 ( .gnd(gnd), .vdd(vdd), .A(_16186_), .B(_16192_), .Y(_16450_) );
	NOR2X1 NOR2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_14564_), .Y(_16451_) );
	NAND2X1 NAND2X1_3268 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_9_bF_buf1), .B(adder_bOperand_22_bF_buf3), .Y(_16452_) );
	NOR2X1 NOR2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_16142_), .B(_16452_), .Y(_16453_) );
	AOI22X1 AOI22X1_373 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf1), .B(adder_bOperand_22_bF_buf2), .C(aOperand_frameOut_9_bF_buf0), .D(adder_bOperand_21_bF_buf2), .Y(_16454_) );
	NOR2X1 NOR2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_16454_), .B(_16453_), .Y(_16455_) );
	XOR2X1 XOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_16455_), .B(_16451_), .Y(_16456_) );
	OAI21X1 OAI21X1_3468 ( .gnd(gnd), .vdd(vdd), .A(_15863_), .B(_16148_), .C(_16421_), .Y(_16457_) );
	NAND2X1 NAND2X1_3269 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_12_bF_buf0), .B(adder_bOperand_19_bF_buf3), .Y(_16458_) );
	OAI21X1 OAI21X1_3469 ( .gnd(gnd), .vdd(vdd), .A(_17236__bF_buf2), .B(_13338_), .C(_16147_), .Y(_16460_) );
	OAI21X1 OAI21X1_3470 ( .gnd(gnd), .vdd(vdd), .A(_16148_), .B(_16458_), .C(_16460_), .Y(_16461_) );
	OAI21X1 OAI21X1_3471 ( .gnd(gnd), .vdd(vdd), .A(_16940_), .B(_13334_), .C(_16461_), .Y(_16462_) );
	NAND2X1 NAND2X1_3270 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf2), .B(adder_bOperand_20_bF_buf1), .Y(_16463_) );
	OR2X2 OR2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_16461_), .B(_16463_), .Y(_16464_) );
	NAND2X1 NAND2X1_3271 ( .gnd(gnd), .vdd(vdd), .A(_16462_), .B(_16464_), .Y(_16465_) );
	XNOR2X1 XNOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_16457_), .B(_16465_), .Y(_16466_) );
	XNOR2X1 XNOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_16466_), .B(_16456_), .Y(_16467_) );
	NAND3X1 NAND3X1_3434 ( .gnd(gnd), .vdd(vdd), .A(_16166_), .B(_16168_), .C(_16172_), .Y(_16468_) );
	OAI21X1 OAI21X1_3472 ( .gnd(gnd), .vdd(vdd), .A(_16160_), .B(_16173_), .C(_16468_), .Y(_16469_) );
	OAI21X1 OAI21X1_3473 ( .gnd(gnd), .vdd(vdd), .A(_15881_), .B(_16162_), .C(_16168_), .Y(_16471_) );
	NAND2X1 NAND2X1_3272 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_15_bF_buf1), .B(adder_bOperand_16_bF_buf0), .Y(_16472_) );
	OAI21X1 OAI21X1_3474 ( .gnd(gnd), .vdd(vdd), .A(_12233_), .B(_12131_), .C(_16161_), .Y(_16473_) );
	OAI21X1 OAI21X1_3475 ( .gnd(gnd), .vdd(vdd), .A(_16162_), .B(_16472_), .C(_16473_), .Y(_16474_) );
	OAI21X1 OAI21X1_3476 ( .gnd(gnd), .vdd(vdd), .A(_11858_), .B(_12566_), .C(_16474_), .Y(_16475_) );
	NAND2X1 NAND2X1_3273 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf4), .B(adder_bOperand_17_bF_buf1), .Y(_16476_) );
	OR2X2 OR2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_16474_), .B(_16476_), .Y(_16477_) );
	NAND2X1 NAND2X1_3274 ( .gnd(gnd), .vdd(vdd), .A(_16475_), .B(_16477_), .Y(_16478_) );
	NAND3X1 NAND3X1_3435 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf3), .B(aOperand_frameOut_15_bF_buf0), .C(_16205_), .Y(_16479_) );
	OAI21X1 OAI21X1_3477 ( .gnd(gnd), .vdd(vdd), .A(_16170_), .B(_16204_), .C(_16479_), .Y(_16480_) );
	XNOR2X1 XNOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_16480_), .B(_16478_), .Y(_16482_) );
	XOR2X1 XOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_16482_), .B(_16471_), .Y(_16483_) );
	XNOR2X1 XNOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_16483_), .B(_16469_), .Y(_16484_) );
	XOR2X1 XOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_16484_), .B(_16467_), .Y(_16485_) );
	NAND2X1 NAND2X1_3275 ( .gnd(gnd), .vdd(vdd), .A(_16227_), .B(_16232_), .Y(_16486_) );
	NAND2X1 NAND2X1_3276 ( .gnd(gnd), .vdd(vdd), .A(_16486_), .B(_16485_), .Y(_16487_) );
	XNOR2X1 XNOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_16484_), .B(_16467_), .Y(_16488_) );
	INVX1 INVX1_2102 ( .gnd(gnd), .vdd(vdd), .A(_16486_), .Y(_16489_) );
	NAND2X1 NAND2X1_3277 ( .gnd(gnd), .vdd(vdd), .A(_16489_), .B(_16488_), .Y(_16490_) );
	NAND3X1 NAND3X1_3436 ( .gnd(gnd), .vdd(vdd), .A(_16450_), .B(_16490_), .C(_16487_), .Y(_16491_) );
	INVX1 INVX1_2103 ( .gnd(gnd), .vdd(vdd), .A(_16450_), .Y(_16493_) );
	NAND2X1 NAND2X1_3278 ( .gnd(gnd), .vdd(vdd), .A(_16486_), .B(_16488_), .Y(_16494_) );
	NAND2X1 NAND2X1_3279 ( .gnd(gnd), .vdd(vdd), .A(_16489_), .B(_16485_), .Y(_16495_) );
	NAND3X1 NAND3X1_3437 ( .gnd(gnd), .vdd(vdd), .A(_16493_), .B(_16494_), .C(_16495_), .Y(_16496_) );
	NAND2X1 NAND2X1_3280 ( .gnd(gnd), .vdd(vdd), .A(_16491_), .B(_16496_), .Y(_16497_) );
	OAI21X1 OAI21X1_3478 ( .gnd(gnd), .vdd(vdd), .A(_16305_), .B(_16307_), .C(_16303_), .Y(_16498_) );
	INVX1 INVX1_2104 ( .gnd(gnd), .vdd(vdd), .A(_16208_), .Y(_16499_) );
	OAI21X1 OAI21X1_3479 ( .gnd(gnd), .vdd(vdd), .A(_16499_), .B(_16217_), .C(_16220_), .Y(_16500_) );
	NOR2X1 NOR2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_12365_), .B(_12461_), .Y(_16501_) );
	NAND2X1 NAND2X1_3281 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_13_bF_buf2), .B(aOperand_frameOut_18_bF_buf2), .Y(_16502_) );
	NOR2X1 NOR2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_16204_), .B(_16502_), .Y(_16504_) );
	AOI22X1 AOI22X1_374 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf1), .B(aOperand_frameOut_18_bF_buf1), .C(adder_bOperand_13_bF_buf1), .D(aOperand_frameOut_17_bF_buf4), .Y(_16505_) );
	NOR2X1 NOR2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_16505_), .B(_16504_), .Y(_16506_) );
	XNOR2X1 XNOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_16506_), .B(_16501_), .Y(_16507_) );
	OAI21X1 OAI21X1_3480 ( .gnd(gnd), .vdd(vdd), .A(_15931_), .B(_16211_), .C(_16216_), .Y(_16508_) );
	NAND2X1 NAND2X1_3282 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_10_bF_buf0), .B(aOperand_frameOut_21_bF_buf0), .Y(_16509_) );
	OAI21X1 OAI21X1_3481 ( .gnd(gnd), .vdd(vdd), .A(_17025__bF_buf3), .B(_13812_), .C(_16210_), .Y(_16510_) );
	OAI21X1 OAI21X1_3482 ( .gnd(gnd), .vdd(vdd), .A(_16211_), .B(_16509_), .C(_16510_), .Y(_16511_) );
	OAI21X1 OAI21X1_3483 ( .gnd(gnd), .vdd(vdd), .A(_17022__bF_buf2), .B(_13224_), .C(_16511_), .Y(_16512_) );
	NAND2X1 NAND2X1_3283 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf2), .B(aOperand_frameOut_19_bF_buf4), .Y(_16513_) );
	OR2X2 OR2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_16511_), .B(_16513_), .Y(_16515_) );
	NAND2X1 NAND2X1_3284 ( .gnd(gnd), .vdd(vdd), .A(_16512_), .B(_16515_), .Y(_16516_) );
	XOR2X1 XOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_16508_), .B(_16516_), .Y(_16517_) );
	XOR2X1 XOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_16517_), .B(_16507_), .Y(_16518_) );
	NAND3X1 NAND3X1_3438 ( .gnd(gnd), .vdd(vdd), .A(_16249_), .B(_16252_), .C(_16256_), .Y(_16519_) );
	OAI21X1 OAI21X1_3484 ( .gnd(gnd), .vdd(vdd), .A(_16243_), .B(_16260_), .C(_16519_), .Y(_16520_) );
	XOR2X1 XOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_16518_), .B(_16520_), .Y(_16521_) );
	OR2X2 OR2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_16521_), .B(_16500_), .Y(_16522_) );
	NAND2X1 NAND2X1_3285 ( .gnd(gnd), .vdd(vdd), .A(_16500_), .B(_16521_), .Y(_16523_) );
	NAND2X1 NAND2X1_3286 ( .gnd(gnd), .vdd(vdd), .A(_16523_), .B(_16522_), .Y(_16524_) );
	INVX1 INVX1_2105 ( .gnd(gnd), .vdd(vdd), .A(_16524_), .Y(_16526_) );
	OAI21X1 OAI21X1_3485 ( .gnd(gnd), .vdd(vdd), .A(_15962_), .B(_16246_), .C(_16252_), .Y(_16527_) );
	NAND2X1 NAND2X1_3287 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_7_bF_buf5), .B(aOperand_frameOut_24_bF_buf0), .Y(_16528_) );
	OAI21X1 OAI21X1_3486 ( .gnd(gnd), .vdd(vdd), .A(_14684__bF_buf2), .B(_14722_), .C(_16245_), .Y(_16529_) );
	OAI21X1 OAI21X1_3487 ( .gnd(gnd), .vdd(vdd), .A(_16246_), .B(_16528_), .C(_16529_), .Y(_16530_) );
	OAI21X1 OAI21X1_3488 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf2), .B(_14125_), .C(_16530_), .Y(_16531_) );
	NAND2X1 NAND2X1_3288 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_8_bF_buf2), .B(aOperand_frameOut_22_bF_buf3), .Y(_16532_) );
	OR2X2 OR2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_16530_), .B(_16532_), .Y(_16533_) );
	NAND2X1 NAND2X1_3289 ( .gnd(gnd), .vdd(vdd), .A(_16531_), .B(_16533_), .Y(_16534_) );
	INVX1 INVX1_2106 ( .gnd(gnd), .vdd(vdd), .A(_16534_), .Y(_16535_) );
	NAND3X1 NAND3X1_3439 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf2), .B(aOperand_frameOut_24_bF_buf3), .C(_16267_), .Y(_16537_) );
	OAI21X1 OAI21X1_3489 ( .gnd(gnd), .vdd(vdd), .A(_16254_), .B(_16266_), .C(_16537_), .Y(_16538_) );
	NOR2X1 NOR2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_16538_), .B(_16535_), .Y(_16539_) );
	AND2X2 AND2X2_409 ( .gnd(gnd), .vdd(vdd), .A(_16535_), .B(_16538_), .Y(_16540_) );
	NOR2X1 NOR2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_16539_), .B(_16540_), .Y(_16541_) );
	NOR2X1 NOR2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_16527_), .B(_16541_), .Y(_16542_) );
	AND2X2 AND2X2_410 ( .gnd(gnd), .vdd(vdd), .A(_16541_), .B(_16527_), .Y(_16543_) );
	NOR2X1 NOR2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_16542_), .B(_16543_), .Y(_16544_) );
	NOR2X1 NOR2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_16279_), .B(_16272_), .Y(_16545_) );
	NOR2X1 NOR2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_16545_), .B(_16287_), .Y(_16546_) );
	NAND2X1 NAND2X1_3290 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf1), .B(aOperand_frameOut_25_bF_buf1), .Y(_16548_) );
	NAND2X1 NAND2X1_3291 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_4_bF_buf4), .B(aOperand_frameOut_27_), .Y(_16549_) );
	NOR2X1 NOR2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_16266_), .B(_16549_), .Y(_16550_) );
	AOI22X1 AOI22X1_375 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf4), .B(aOperand_frameOut_27_), .C(adder_bOperand_4_bF_buf3), .D(aOperand_frameOut_26_), .Y(_16551_) );
	OAI21X1 OAI21X1_3490 ( .gnd(gnd), .vdd(vdd), .A(_16551_), .B(_16550_), .C(_16548_), .Y(_16552_) );
	NOR2X1 NOR2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_16551_), .B(_16550_), .Y(_16553_) );
	NAND3X1 NAND3X1_3440 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_5_bF_buf0), .B(aOperand_frameOut_25_bF_buf0), .C(_16553_), .Y(_16554_) );
	NAND2X1 NAND2X1_3292 ( .gnd(gnd), .vdd(vdd), .A(_16552_), .B(_16554_), .Y(_16555_) );
	OAI22X1 OAI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_16269_), .B(_16275_), .C(_16274_), .D(_16278_), .Y(_16556_) );
	NAND2X1 NAND2X1_3293 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf4), .B(aOperand_frameOut_28_), .Y(_16557_) );
	NAND2X1 NAND2X1_3294 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_1_bF_buf4), .B(aOperand_frameOut_30_), .Y(_16559_) );
	INVX1 INVX1_2107 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_30_), .Y(_16560_) );
	OAI21X1 OAI21X1_3491 ( .gnd(gnd), .vdd(vdd), .A(_17295__bF_buf0), .B(_16560_), .C(_16275_), .Y(_16561_) );
	OAI21X1 OAI21X1_3492 ( .gnd(gnd), .vdd(vdd), .A(_16276_), .B(_16559_), .C(_16561_), .Y(_16562_) );
	XOR2X1 XOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_16562_), .B(_16557_), .Y(_16563_) );
	XNOR2X1 XNOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_16563_), .B(_16556_), .Y(_16564_) );
	XNOR2X1 XNOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_16564_), .B(_16555_), .Y(_16565_) );
	OR2X2 OR2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_16546_), .B(_16565_), .Y(_16566_) );
	NAND2X1 NAND2X1_3295 ( .gnd(gnd), .vdd(vdd), .A(_16565_), .B(_16546_), .Y(_16567_) );
	NAND3X1 NAND3X1_3441 ( .gnd(gnd), .vdd(vdd), .A(_16567_), .B(_16566_), .C(_16544_), .Y(_16568_) );
	NAND2X1 NAND2X1_3296 ( .gnd(gnd), .vdd(vdd), .A(_16567_), .B(_16566_), .Y(_16570_) );
	OAI21X1 OAI21X1_3493 ( .gnd(gnd), .vdd(vdd), .A(_16542_), .B(_16543_), .C(_16570_), .Y(_16571_) );
	AND2X2 AND2X2_411 ( .gnd(gnd), .vdd(vdd), .A(_16571_), .B(_16568_), .Y(_16572_) );
	OAI21X1 OAI21X1_3494 ( .gnd(gnd), .vdd(vdd), .A(_16297_), .B(_16298_), .C(_16572_), .Y(_16573_) );
	OAI21X1 OAI21X1_3495 ( .gnd(gnd), .vdd(vdd), .A(_16294_), .B(_16296_), .C(_16292_), .Y(_16574_) );
	INVX1 INVX1_2108 ( .gnd(gnd), .vdd(vdd), .A(_16574_), .Y(_16575_) );
	NAND2X1 NAND2X1_3297 ( .gnd(gnd), .vdd(vdd), .A(_16568_), .B(_16571_), .Y(_16576_) );
	NAND2X1 NAND2X1_3298 ( .gnd(gnd), .vdd(vdd), .A(_16575_), .B(_16576_), .Y(_16577_) );
	NAND3X1 NAND3X1_3442 ( .gnd(gnd), .vdd(vdd), .A(_16573_), .B(_16577_), .C(_16526_), .Y(_16578_) );
	NOR2X1 NOR2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_16575_), .B(_16576_), .Y(_16579_) );
	NOR2X1 NOR2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_16574_), .B(_16572_), .Y(_16581_) );
	OAI21X1 OAI21X1_3496 ( .gnd(gnd), .vdd(vdd), .A(_16579_), .B(_16581_), .C(_16524_), .Y(_16582_) );
	NAND3X1 NAND3X1_3443 ( .gnd(gnd), .vdd(vdd), .A(_16498_), .B(_16578_), .C(_16582_), .Y(_16583_) );
	INVX1 INVX1_2109 ( .gnd(gnd), .vdd(vdd), .A(_16498_), .Y(_16584_) );
	NAND2X1 NAND2X1_3299 ( .gnd(gnd), .vdd(vdd), .A(_16575_), .B(_16572_), .Y(_16585_) );
	OAI21X1 OAI21X1_3497 ( .gnd(gnd), .vdd(vdd), .A(_16297_), .B(_16298_), .C(_16576_), .Y(_16586_) );
	AOI21X1 AOI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_16585_), .B(_16586_), .C(_16524_), .Y(_16587_) );
	AOI21X1 AOI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_16573_), .B(_16577_), .C(_16526_), .Y(_16588_) );
	OAI21X1 OAI21X1_3498 ( .gnd(gnd), .vdd(vdd), .A(_16587_), .B(_16588_), .C(_16584_), .Y(_16589_) );
	NAND3X1 NAND3X1_3444 ( .gnd(gnd), .vdd(vdd), .A(_16497_), .B(_16583_), .C(_16589_), .Y(_16590_) );
	AND2X2 AND2X2_412 ( .gnd(gnd), .vdd(vdd), .A(_16491_), .B(_16496_), .Y(_16592_) );
	NAND3X1 NAND3X1_3445 ( .gnd(gnd), .vdd(vdd), .A(_16584_), .B(_16578_), .C(_16582_), .Y(_16593_) );
	OAI21X1 OAI21X1_3499 ( .gnd(gnd), .vdd(vdd), .A(_16587_), .B(_16588_), .C(_16498_), .Y(_16594_) );
	NAND3X1 NAND3X1_3446 ( .gnd(gnd), .vdd(vdd), .A(_16593_), .B(_16592_), .C(_16594_), .Y(_16595_) );
	NAND2X1 NAND2X1_3300 ( .gnd(gnd), .vdd(vdd), .A(_16590_), .B(_16595_), .Y(_16596_) );
	OAI21X1 OAI21X1_3500 ( .gnd(gnd), .vdd(vdd), .A(_16319_), .B(_16320_), .C(_16596_), .Y(_16597_) );
	OAI21X1 OAI21X1_3501 ( .gnd(gnd), .vdd(vdd), .A(_16318_), .B(_16316_), .C(_16314_), .Y(_16598_) );
	INVX1 INVX1_2110 ( .gnd(gnd), .vdd(vdd), .A(_16598_), .Y(_16599_) );
	NAND3X1 NAND3X1_3447 ( .gnd(gnd), .vdd(vdd), .A(_16583_), .B(_16592_), .C(_16589_), .Y(_16600_) );
	NAND3X1 NAND3X1_3448 ( .gnd(gnd), .vdd(vdd), .A(_16497_), .B(_16593_), .C(_16594_), .Y(_16601_) );
	NAND2X1 NAND2X1_3301 ( .gnd(gnd), .vdd(vdd), .A(_16601_), .B(_16600_), .Y(_16603_) );
	NAND2X1 NAND2X1_3302 ( .gnd(gnd), .vdd(vdd), .A(_16599_), .B(_16603_), .Y(_16604_) );
	NAND3X1 NAND3X1_3449 ( .gnd(gnd), .vdd(vdd), .A(_16449_), .B(_16604_), .C(_16597_), .Y(_16605_) );
	NAND3X1 NAND3X1_3450 ( .gnd(gnd), .vdd(vdd), .A(_16444_), .B(_16438_), .C(_16442_), .Y(_16606_) );
	NAND3X1 NAND3X1_3451 ( .gnd(gnd), .vdd(vdd), .A(_16381_), .B(_16446_), .C(_16445_), .Y(_16607_) );
	NAND2X1 NAND2X1_3303 ( .gnd(gnd), .vdd(vdd), .A(_16606_), .B(_16607_), .Y(_16608_) );
	NAND2X1 NAND2X1_3304 ( .gnd(gnd), .vdd(vdd), .A(_16599_), .B(_16596_), .Y(_16609_) );
	OAI21X1 OAI21X1_3502 ( .gnd(gnd), .vdd(vdd), .A(_16319_), .B(_16320_), .C(_16603_), .Y(_16610_) );
	NAND3X1 NAND3X1_3452 ( .gnd(gnd), .vdd(vdd), .A(_16608_), .B(_16609_), .C(_16610_), .Y(_16611_) );
	NAND2X1 NAND2X1_3305 ( .gnd(gnd), .vdd(vdd), .A(_16605_), .B(_16611_), .Y(_16612_) );
	NAND2X1 NAND2X1_3306 ( .gnd(gnd), .vdd(vdd), .A(_16380_), .B(_16612_), .Y(_16614_) );
	AOI21X1 AOI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_16610_), .B(_16609_), .C(_16449_), .Y(_16615_) );
	AOI21X1 AOI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_16597_), .B(_16604_), .C(_16608_), .Y(_16616_) );
	OAI21X1 OAI21X1_3503 ( .gnd(gnd), .vdd(vdd), .A(_16616_), .B(_16615_), .C(_16379_), .Y(_16617_) );
	AOI21X1 AOI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_16614_), .B(_16617_), .C(_16378_), .Y(_16618_) );
	AOI21X1 AOI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_16605_), .B(_16611_), .C(_16380_), .Y(_16619_) );
	NAND3X1 NAND3X1_3453 ( .gnd(gnd), .vdd(vdd), .A(_16608_), .B(_16604_), .C(_16597_), .Y(_16620_) );
	NAND3X1 NAND3X1_3454 ( .gnd(gnd), .vdd(vdd), .A(_16449_), .B(_16609_), .C(_16610_), .Y(_16621_) );
	AOI21X1 AOI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_16621_), .B(_16620_), .C(_16379_), .Y(_16622_) );
	OAI21X1 OAI21X1_3504 ( .gnd(gnd), .vdd(vdd), .A(_16619_), .B(_16622_), .C(_16378_), .Y(_16623_) );
	INVX1 INVX1_2111 ( .gnd(gnd), .vdd(vdd), .A(_16623_), .Y(_16625_) );
	OAI21X1 OAI21X1_3505 ( .gnd(gnd), .vdd(vdd), .A(_16618_), .B(_16625_), .C(_16377_), .Y(_16626_) );
	INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(_16377_), .Y(_16627_) );
	INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(_16378_), .Y(_16628_) );
	AOI21X1 AOI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_16614_), .B(_16617_), .C(_16628_), .Y(_16629_) );
	NAND2X1 NAND2X1_3307 ( .gnd(gnd), .vdd(vdd), .A(_16379_), .B(_16612_), .Y(_16630_) );
	OAI21X1 OAI21X1_3506 ( .gnd(gnd), .vdd(vdd), .A(_16615_), .B(_16616_), .C(_16380_), .Y(_16631_) );
	AOI21X1 AOI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_16630_), .B(_16631_), .C(_16378_), .Y(_16632_) );
	OAI21X1 OAI21X1_3507 ( .gnd(gnd), .vdd(vdd), .A(_16629_), .B(_16632_), .C(_16627_), .Y(_16633_) );
	NAND3X1 NAND3X1_3455 ( .gnd(gnd), .vdd(vdd), .A(_16343_), .B(_16633_), .C(_16626_), .Y(_16634_) );
	INVX1 INVX1_2112 ( .gnd(gnd), .vdd(vdd), .A(_16343_), .Y(_16636_) );
	OAI21X1 OAI21X1_3508 ( .gnd(gnd), .vdd(vdd), .A(_16618_), .B(_16625_), .C(_16627_), .Y(_16637_) );
	OAI21X1 OAI21X1_3509 ( .gnd(gnd), .vdd(vdd), .A(_16629_), .B(_16632_), .C(_16377_), .Y(_16638_) );
	NAND3X1 NAND3X1_3456 ( .gnd(gnd), .vdd(vdd), .A(_16636_), .B(_16638_), .C(_16637_), .Y(_16639_) );
	AOI22X1 AOI22X1_376 ( .gnd(gnd), .vdd(vdd), .A(_16634_), .B(_16639_), .C(_16376_), .D(_16374_), .Y(_16640_) );
	NAND2X1 NAND2X1_3308 ( .gnd(gnd), .vdd(vdd), .A(_16376_), .B(_16374_), .Y(_16641_) );
	NAND2X1 NAND2X1_3309 ( .gnd(gnd), .vdd(vdd), .A(_16634_), .B(_16639_), .Y(_16642_) );
	NOR2X1 NOR2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_16642_), .B(_16641_), .Y(_16643_) );
	NOR2X1 NOR2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_16640_), .B(_16643_), .Y(mulOut_30_) );
	NAND2X1 NAND2X1_3310 ( .gnd(gnd), .vdd(vdd), .A(_16633_), .B(_16626_), .Y(_16644_) );
	NOR2X1 NOR2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_16343_), .B(_16644_), .Y(_16646_) );
	INVX1 INVX1_2113 ( .gnd(gnd), .vdd(vdd), .A(_16646_), .Y(_16647_) );
	NOR2X1 NOR2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_15126_), .B(_15784_), .Y(_16648_) );
	OAI21X1 OAI21X1_3510 ( .gnd(gnd), .vdd(vdd), .A(_14538_), .B(_14532_), .C(_16648_), .Y(_16649_) );
	AND2X2 AND2X2_413 ( .gnd(gnd), .vdd(vdd), .A(_16060_), .B(_16063_), .Y(_16650_) );
	NAND2X1 NAND2X1_3311 ( .gnd(gnd), .vdd(vdd), .A(_16355_), .B(_16650_), .Y(_16651_) );
	AOI21X1 AOI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_16649_), .B(_15787_), .C(_16651_), .Y(_16652_) );
	INVX1 INVX1_2114 ( .gnd(gnd), .vdd(vdd), .A(_16375_), .Y(_16653_) );
	NAND2X1 NAND2X1_3312 ( .gnd(gnd), .vdd(vdd), .A(_16066_), .B(_16355_), .Y(_16654_) );
	NAND2X1 NAND2X1_3313 ( .gnd(gnd), .vdd(vdd), .A(_16653_), .B(_16654_), .Y(_16655_) );
	OAI21X1 OAI21X1_3511 ( .gnd(gnd), .vdd(vdd), .A(_16655_), .B(_16652_), .C(_16642_), .Y(_16657_) );
	OAI21X1 OAI21X1_3512 ( .gnd(gnd), .vdd(vdd), .A(_16628_), .B(_16622_), .C(_16630_), .Y(_16658_) );
	NAND2X1 NAND2X1_3314 ( .gnd(gnd), .vdd(vdd), .A(_16438_), .B(_16443_), .Y(_16659_) );
	INVX1 INVX1_2115 ( .gnd(gnd), .vdd(vdd), .A(_16659_), .Y(_16660_) );
	NOR2X1 NOR2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_16598_), .B(_16596_), .Y(_16661_) );
	OAI21X1 OAI21X1_3513 ( .gnd(gnd), .vdd(vdd), .A(_16449_), .B(_16661_), .C(_16597_), .Y(_16662_) );
	NOR2X1 NOR2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_16489_), .B(_16488_), .Y(_16663_) );
	AOI21X1 AOI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_16450_), .B(_16490_), .C(_16663_), .Y(_16664_) );
	OAI21X1 OAI21X1_3514 ( .gnd(gnd), .vdd(vdd), .A(_16076_), .B(_16388_), .C(_16392_), .Y(_16665_) );
	NAND2X1 NAND2X1_3315 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_4_bF_buf3), .B(adder_bOperand_27_), .Y(_16666_) );
	XNOR2X1 XNOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_16388_), .B(_16666_), .Y(_16668_) );
	NAND2X1 NAND2X1_3316 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_1_bF_buf0), .B(adder_bOperand_30_), .Y(_16669_) );
	NAND2X1 NAND2X1_3317 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_2_bF_buf4), .B(adder_bOperand_29_), .Y(_16670_) );
	XNOR2X1 XNOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_16669_), .B(_16670_), .Y(_16671_) );
	XNOR2X1 XNOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_16668_), .B(_16671_), .Y(_16672_) );
	XNOR2X1 XNOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_16672_), .B(_16665_), .Y(_16673_) );
	OAI21X1 OAI21X1_3515 ( .gnd(gnd), .vdd(vdd), .A(_16383_), .B(_16396_), .C(_16394_), .Y(_16674_) );
	XNOR2X1 XNOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_16674_), .B(_16673_), .Y(_16675_) );
	NAND3X1 NAND3X1_3457 ( .gnd(gnd), .vdd(vdd), .A(_16462_), .B(_16464_), .C(_16457_), .Y(_16676_) );
	NAND2X1 NAND2X1_3318 ( .gnd(gnd), .vdd(vdd), .A(_16456_), .B(_16466_), .Y(_16677_) );
	OAI22X1 OAI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(_16089_), .B(_16410_), .C(_16409_), .D(_16412_), .Y(_16679_) );
	AOI21X1 AOI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_16455_), .B(_16451_), .C(_16453_), .Y(_16680_) );
	NOR2X1 NOR2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_12780_), .B(_15806_), .Y(_16681_) );
	NAND2X1 NAND2X1_3319 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_7_bF_buf1), .B(adder_bOperand_24_), .Y(_16682_) );
	XNOR2X1 XNOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_16410_), .B(_16682_), .Y(_16683_) );
	XNOR2X1 XNOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_16683_), .B(_16681_), .Y(_16684_) );
	XOR2X1 XOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_16684_), .B(_16680_), .Y(_16685_) );
	XNOR2X1 XNOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_16685_), .B(_16679_), .Y(_16686_) );
	NAND3X1 NAND3X1_3458 ( .gnd(gnd), .vdd(vdd), .A(_16676_), .B(_16677_), .C(_16686_), .Y(_16687_) );
	NAND2X1 NAND2X1_3320 ( .gnd(gnd), .vdd(vdd), .A(_16676_), .B(_16677_), .Y(_16688_) );
	XOR2X1 XOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_16685_), .B(_16679_), .Y(_16690_) );
	NAND2X1 NAND2X1_3321 ( .gnd(gnd), .vdd(vdd), .A(_16690_), .B(_16688_), .Y(_16691_) );
	NAND2X1 NAND2X1_3322 ( .gnd(gnd), .vdd(vdd), .A(_16691_), .B(_16687_), .Y(_16692_) );
	INVX1 INVX1_2116 ( .gnd(gnd), .vdd(vdd), .A(_16413_), .Y(_16693_) );
	NAND2X1 NAND2X1_3323 ( .gnd(gnd), .vdd(vdd), .A(_16417_), .B(_16693_), .Y(_16694_) );
	NAND2X1 NAND2X1_3324 ( .gnd(gnd), .vdd(vdd), .A(_16408_), .B(_16418_), .Y(_16695_) );
	NAND2X1 NAND2X1_3325 ( .gnd(gnd), .vdd(vdd), .A(_16694_), .B(_16695_), .Y(_16696_) );
	XOR2X1 XOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_16692_), .B(_16696_), .Y(_16697_) );
	XNOR2X1 XNOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_16697_), .B(_16675_), .Y(_16698_) );
	NAND2X1 NAND2X1_3326 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_0_bF_buf2), .B(divider_absoluteValue_B_msb), .Y(_16699_) );
	OAI21X1 OAI21X1_3516 ( .gnd(gnd), .vdd(vdd), .A(_16407_), .B(_16425_), .C(_16430_), .Y(_16701_) );
	XOR2X1 XOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_16701_), .B(_16699_), .Y(_16702_) );
	NAND2X1 NAND2X1_3327 ( .gnd(gnd), .vdd(vdd), .A(_16702_), .B(_16698_), .Y(_16703_) );
	XOR2X1 XOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_16697_), .B(_16675_), .Y(_16704_) );
	XNOR2X1 XNOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_16701_), .B(_16699_), .Y(_16705_) );
	NAND2X1 NAND2X1_3328 ( .gnd(gnd), .vdd(vdd), .A(_16705_), .B(_16704_), .Y(_16706_) );
	NAND3X1 NAND3X1_3459 ( .gnd(gnd), .vdd(vdd), .A(_16664_), .B(_16703_), .C(_16706_), .Y(_16707_) );
	INVX1 INVX1_2117 ( .gnd(gnd), .vdd(vdd), .A(_16664_), .Y(_16708_) );
	NAND2X1 NAND2X1_3329 ( .gnd(gnd), .vdd(vdd), .A(_16702_), .B(_16704_), .Y(_16709_) );
	NAND2X1 NAND2X1_3330 ( .gnd(gnd), .vdd(vdd), .A(_16705_), .B(_16698_), .Y(_16710_) );
	NAND3X1 NAND3X1_3460 ( .gnd(gnd), .vdd(vdd), .A(_16710_), .B(_16709_), .C(_16708_), .Y(_16712_) );
	INVX1 INVX1_2118 ( .gnd(gnd), .vdd(vdd), .A(_16402_), .Y(_16713_) );
	NOR2X1 NOR2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_16432_), .B(_16713_), .Y(_16714_) );
	INVX1 INVX1_2119 ( .gnd(gnd), .vdd(vdd), .A(_16714_), .Y(_16715_) );
	OAI21X1 OAI21X1_3517 ( .gnd(gnd), .vdd(vdd), .A(_16401_), .B(_16433_), .C(_16715_), .Y(_16716_) );
	NAND3X1 NAND3X1_3461 ( .gnd(gnd), .vdd(vdd), .A(_16716_), .B(_16707_), .C(_16712_), .Y(_16717_) );
	NAND3X1 NAND3X1_3462 ( .gnd(gnd), .vdd(vdd), .A(_16664_), .B(_16710_), .C(_16709_), .Y(_16718_) );
	NAND3X1 NAND3X1_3463 ( .gnd(gnd), .vdd(vdd), .A(_16706_), .B(_16703_), .C(_16708_), .Y(_16719_) );
	INVX1 INVX1_2120 ( .gnd(gnd), .vdd(vdd), .A(_16716_), .Y(_16720_) );
	NAND3X1 NAND3X1_3464 ( .gnd(gnd), .vdd(vdd), .A(_16718_), .B(_16720_), .C(_16719_), .Y(_16721_) );
	AND2X2 AND2X2_414 ( .gnd(gnd), .vdd(vdd), .A(_16721_), .B(_16717_), .Y(_16723_) );
	NAND2X1 NAND2X1_3331 ( .gnd(gnd), .vdd(vdd), .A(_16469_), .B(_16483_), .Y(_16724_) );
	OAI21X1 OAI21X1_3518 ( .gnd(gnd), .vdd(vdd), .A(_16467_), .B(_16484_), .C(_16724_), .Y(_16725_) );
	NAND2X1 NAND2X1_3332 ( .gnd(gnd), .vdd(vdd), .A(_16520_), .B(_16518_), .Y(_16726_) );
	NAND2X1 NAND2X1_3333 ( .gnd(gnd), .vdd(vdd), .A(_16726_), .B(_16523_), .Y(_16727_) );
	AOI21X1 AOI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_16506_), .B(_16501_), .C(_16504_), .Y(_16728_) );
	NAND2X1 NAND2X1_3334 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_14_bF_buf0), .B(adder_bOperand_17_bF_buf0), .Y(_16729_) );
	NAND2X1 NAND2X1_3335 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_15_bF_buf0), .B(aOperand_frameOut_16_bF_buf0), .Y(_16730_) );
	XNOR2X1 XNOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_16472_), .B(_16730_), .Y(_16731_) );
	XNOR2X1 XNOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_16731_), .B(_16729_), .Y(_16732_) );
	XOR2X1 XOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_16732_), .B(_16728_), .Y(_16734_) );
	NAND2X1 NAND2X1_3336 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_10_bF_buf1), .B(adder_bOperand_21_bF_buf1), .Y(_16735_) );
	XNOR2X1 XNOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_16452_), .B(_16735_), .Y(_16736_) );
	NAND2X1 NAND2X1_3337 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_11_bF_buf0), .B(adder_bOperand_20_bF_buf0), .Y(_16737_) );
	NAND2X1 NAND2X1_3338 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_13_bF_buf3), .B(adder_bOperand_18_bF_buf3), .Y(_16738_) );
	XNOR2X1 XNOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_16458_), .B(_16738_), .Y(_16739_) );
	XNOR2X1 XNOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_16739_), .B(_16737_), .Y(_16740_) );
	XNOR2X1 XNOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_16740_), .B(_16736_), .Y(_16741_) );
	OAI21X1 OAI21X1_3519 ( .gnd(gnd), .vdd(vdd), .A(_16162_), .B(_16472_), .C(_16477_), .Y(_16742_) );
	XNOR2X1 XNOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_16741_), .B(_16742_), .Y(_16743_) );
	XNOR2X1 XNOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_16743_), .B(_16734_), .Y(_16745_) );
	NAND2X1 NAND2X1_3339 ( .gnd(gnd), .vdd(vdd), .A(aOperand_frameOut_8_bF_buf0), .B(adder_bOperand_23_), .Y(_16746_) );
	OAI21X1 OAI21X1_3520 ( .gnd(gnd), .vdd(vdd), .A(_16148_), .B(_16458_), .C(_16464_), .Y(_16747_) );
	XNOR2X1 XNOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_16747_), .B(_16746_), .Y(_16748_) );
	NAND3X1 NAND3X1_3465 ( .gnd(gnd), .vdd(vdd), .A(_16475_), .B(_16477_), .C(_16480_), .Y(_16749_) );
	NAND2X1 NAND2X1_3340 ( .gnd(gnd), .vdd(vdd), .A(_16471_), .B(_16482_), .Y(_16750_) );
	NAND2X1 NAND2X1_3341 ( .gnd(gnd), .vdd(vdd), .A(_16749_), .B(_16750_), .Y(_16751_) );
	XNOR2X1 XNOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_16751_), .B(_16748_), .Y(_16752_) );
	XNOR2X1 XNOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_16752_), .B(_16745_), .Y(_16753_) );
	NOR2X1 NOR2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_16727_), .B(_16753_), .Y(_16754_) );
	NAND2X1 NAND2X1_3342 ( .gnd(gnd), .vdd(vdd), .A(_16727_), .B(_16753_), .Y(_16756_) );
	INVX1 INVX1_2121 ( .gnd(gnd), .vdd(vdd), .A(_16756_), .Y(_16757_) );
	OAI21X1 OAI21X1_3521 ( .gnd(gnd), .vdd(vdd), .A(_16754_), .B(_16757_), .C(_16725_), .Y(_16758_) );
	INVX1 INVX1_2122 ( .gnd(gnd), .vdd(vdd), .A(_16725_), .Y(_16759_) );
	INVX1 INVX1_2123 ( .gnd(gnd), .vdd(vdd), .A(_16754_), .Y(_16760_) );
	NAND3X1 NAND3X1_3466 ( .gnd(gnd), .vdd(vdd), .A(_16759_), .B(_16756_), .C(_16760_), .Y(_16761_) );
	AND2X2 AND2X2_415 ( .gnd(gnd), .vdd(vdd), .A(_16761_), .B(_16758_), .Y(_16762_) );
	AOI21X1 AOI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_16526_), .B(_16577_), .C(_16579_), .Y(_16763_) );
	INVX1 INVX1_2124 ( .gnd(gnd), .vdd(vdd), .A(_16516_), .Y(_16764_) );
	NOR2X1 NOR2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_16507_), .B(_16517_), .Y(_16765_) );
	AOI21X1 AOI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_16508_), .B(_16764_), .C(_16765_), .Y(_16767_) );
	NAND2X1 NAND2X1_3343 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_12_bF_buf0), .B(aOperand_frameOut_19_bF_buf3), .Y(_16768_) );
	XOR2X1 XOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_16502_), .B(_16768_), .Y(_16769_) );
	NAND2X1 NAND2X1_3344 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_11_bF_buf1), .B(aOperand_frameOut_20_bF_buf0), .Y(_16770_) );
	NAND2X1 NAND2X1_3345 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_9_bF_buf2), .B(aOperand_frameOut_22_bF_buf2), .Y(_16771_) );
	XNOR2X1 XNOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_16509_), .B(_16771_), .Y(_16772_) );
	XNOR2X1 XNOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_16772_), .B(_16770_), .Y(_16773_) );
	XNOR2X1 XNOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_16773_), .B(_16769_), .Y(_16774_) );
	NAND2X1 NAND2X1_3346 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_14_bF_buf2), .B(aOperand_frameOut_17_bF_buf3), .Y(_16775_) );
	OAI21X1 OAI21X1_3522 ( .gnd(gnd), .vdd(vdd), .A(_16211_), .B(_16509_), .C(_16515_), .Y(_16776_) );
	XNOR2X1 XNOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_16776_), .B(_16775_), .Y(_16778_) );
	XNOR2X1 XNOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_16778_), .B(_16774_), .Y(_16779_) );
	OR2X2 OR2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_16543_), .B(_16540_), .Y(_16780_) );
	XNOR2X1 XNOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_16780_), .B(_16779_), .Y(_16781_) );
	XNOR2X1 XNOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_16781_), .B(_16767_), .Y(_16782_) );
	OAI21X1 OAI21X1_3523 ( .gnd(gnd), .vdd(vdd), .A(_16546_), .B(_16565_), .C(_16568_), .Y(_16783_) );
	OAI21X1 OAI21X1_3524 ( .gnd(gnd), .vdd(vdd), .A(_16266_), .B(_16549_), .C(_16554_), .Y(_16784_) );
	NOR2X1 NOR2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_14728__bF_buf1), .B(_14436_), .Y(_16785_) );
	NAND2X1 NAND2X1_3347 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_6_bF_buf5), .B(aOperand_frameOut_25_bF_buf3), .Y(_16786_) );
	XNOR2X1 XNOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_16528_), .B(_16786_), .Y(_16787_) );
	XNOR2X1 XNOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_16787_), .B(_16785_), .Y(_16789_) );
	XNOR2X1 XNOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_16789_), .B(_16784_), .Y(_16790_) );
	NOR2X1 NOR2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_13436__bF_buf2), .B(_15674_), .Y(_16791_) );
	NAND2X1 NAND2X1_3348 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_3_bF_buf3), .B(aOperand_frameOut_28_), .Y(_16792_) );
	XNOR2X1 XNOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_16549_), .B(_16792_), .Y(_16793_) );
	XNOR2X1 XNOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_16793_), .B(_16791_), .Y(_16794_) );
	OAI22X1 OAI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_16276_), .B(_16559_), .C(_16557_), .D(_16562_), .Y(_16795_) );
	NAND2X1 NAND2X1_3349 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_2_bF_buf3), .B(aOperand_frameOut_29_), .Y(_16796_) );
	NAND2X1 NAND2X1_3350 ( .gnd(gnd), .vdd(vdd), .A(adder_bOperand_0_bF_buf1), .B(divider_absoluteValue_A_msb), .Y(_16797_) );
	XNOR2X1 XNOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_16559_), .B(_16797_), .Y(_16798_) );
	XNOR2X1 XNOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_16798_), .B(_16796_), .Y(_16800_) );
	XNOR2X1 XNOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_16800_), .B(_16795_), .Y(_16801_) );
	XNOR2X1 XNOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_16801_), .B(_16794_), .Y(_16802_) );
	XNOR2X1 XNOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_16802_), .B(_16790_), .Y(_16803_) );
	OAI21X1 OAI21X1_3525 ( .gnd(gnd), .vdd(vdd), .A(_16246_), .B(_16528_), .C(_16533_), .Y(_16804_) );
	NAND2X1 NAND2X1_3351 ( .gnd(gnd), .vdd(vdd), .A(_16556_), .B(_16563_), .Y(_16805_) );
	OAI21X1 OAI21X1_3526 ( .gnd(gnd), .vdd(vdd), .A(_16555_), .B(_16564_), .C(_16805_), .Y(_16806_) );
	XNOR2X1 XNOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_16806_), .B(_16804_), .Y(_16807_) );
	XOR2X1 XOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_16803_), .B(_16807_), .Y(_16808_) );
	NAND2X1 NAND2X1_3352 ( .gnd(gnd), .vdd(vdd), .A(_16783_), .B(_16808_), .Y(_16809_) );
	INVX1 INVX1_2125 ( .gnd(gnd), .vdd(vdd), .A(_16809_), .Y(_16811_) );
	NOR2X1 NOR2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_16783_), .B(_16808_), .Y(_16812_) );
	OAI21X1 OAI21X1_3527 ( .gnd(gnd), .vdd(vdd), .A(_16812_), .B(_16811_), .C(_16782_), .Y(_16813_) );
	XOR2X1 XOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_16781_), .B(_16767_), .Y(_16814_) );
	INVX1 INVX1_2126 ( .gnd(gnd), .vdd(vdd), .A(_16812_), .Y(_16815_) );
	NAND3X1 NAND3X1_3467 ( .gnd(gnd), .vdd(vdd), .A(_16814_), .B(_16809_), .C(_16815_), .Y(_16816_) );
	AOI21X1 AOI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_16816_), .B(_16813_), .C(_16763_), .Y(_16817_) );
	OAI21X1 OAI21X1_3528 ( .gnd(gnd), .vdd(vdd), .A(_16524_), .B(_16581_), .C(_16573_), .Y(_16818_) );
	XNOR2X1 XNOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_16783_), .B(_16767_), .Y(_16819_) );
	NAND2X1 NAND2X1_3353 ( .gnd(gnd), .vdd(vdd), .A(_16781_), .B(_16808_), .Y(_16820_) );
	INVX1 INVX1_2127 ( .gnd(gnd), .vdd(vdd), .A(_16781_), .Y(_16822_) );
	XNOR2X1 XNOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_16803_), .B(_16807_), .Y(_16823_) );
	NAND2X1 NAND2X1_3354 ( .gnd(gnd), .vdd(vdd), .A(_16823_), .B(_16822_), .Y(_16824_) );
	NAND3X1 NAND3X1_3468 ( .gnd(gnd), .vdd(vdd), .A(_16820_), .B(_16824_), .C(_16819_), .Y(_16825_) );
	INVX1 INVX1_2128 ( .gnd(gnd), .vdd(vdd), .A(_16819_), .Y(_16826_) );
	NAND2X1 NAND2X1_3355 ( .gnd(gnd), .vdd(vdd), .A(_16820_), .B(_16824_), .Y(_16827_) );
	NAND2X1 NAND2X1_3356 ( .gnd(gnd), .vdd(vdd), .A(_16826_), .B(_16827_), .Y(_16828_) );
	AOI21X1 AOI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_16828_), .B(_16825_), .C(_16818_), .Y(_16829_) );
	OAI21X1 OAI21X1_3529 ( .gnd(gnd), .vdd(vdd), .A(_16817_), .B(_16829_), .C(_16762_), .Y(_16830_) );
	NAND2X1 NAND2X1_3357 ( .gnd(gnd), .vdd(vdd), .A(_16758_), .B(_16761_), .Y(_16831_) );
	NAND3X1 NAND3X1_3469 ( .gnd(gnd), .vdd(vdd), .A(_16818_), .B(_16825_), .C(_16828_), .Y(_16833_) );
	NAND3X1 NAND3X1_3470 ( .gnd(gnd), .vdd(vdd), .A(_16763_), .B(_16813_), .C(_16816_), .Y(_16834_) );
	NAND3X1 NAND3X1_3471 ( .gnd(gnd), .vdd(vdd), .A(_16834_), .B(_16833_), .C(_16831_), .Y(_16835_) );
	AOI22X1 AOI22X1_377 ( .gnd(gnd), .vdd(vdd), .A(_16583_), .B(_16600_), .C(_16835_), .D(_16830_), .Y(_16836_) );
	XNOR2X1 XNOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_16818_), .B(_16759_), .Y(_16837_) );
	NAND2X1 NAND2X1_3358 ( .gnd(gnd), .vdd(vdd), .A(_16756_), .B(_16760_), .Y(_16838_) );
	NAND3X1 NAND3X1_3472 ( .gnd(gnd), .vdd(vdd), .A(_16825_), .B(_16828_), .C(_16838_), .Y(_16839_) );
	NOR2X1 NOR2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_16754_), .B(_16757_), .Y(_16840_) );
	NAND3X1 NAND3X1_3473 ( .gnd(gnd), .vdd(vdd), .A(_16813_), .B(_16816_), .C(_16840_), .Y(_16841_) );
	NAND3X1 NAND3X1_3474 ( .gnd(gnd), .vdd(vdd), .A(_16839_), .B(_16841_), .C(_16837_), .Y(_16842_) );
	XNOR2X1 XNOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_16818_), .B(_16725_), .Y(_16844_) );
	AOI21X1 AOI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_16816_), .B(_16813_), .C(_16840_), .Y(_16845_) );
	AOI21X1 AOI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_16828_), .B(_16825_), .C(_16838_), .Y(_16846_) );
	OAI21X1 OAI21X1_3530 ( .gnd(gnd), .vdd(vdd), .A(_16845_), .B(_16846_), .C(_16844_), .Y(_16847_) );
	NAND2X1 NAND2X1_3359 ( .gnd(gnd), .vdd(vdd), .A(_16583_), .B(_16600_), .Y(_16848_) );
	AOI21X1 AOI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_16842_), .B(_16847_), .C(_16848_), .Y(_16849_) );
	OAI21X1 OAI21X1_3531 ( .gnd(gnd), .vdd(vdd), .A(_16836_), .B(_16849_), .C(_16723_), .Y(_16850_) );
	INVX1 INVX1_2129 ( .gnd(gnd), .vdd(vdd), .A(_16723_), .Y(_16851_) );
	NAND3X1 NAND3X1_3475 ( .gnd(gnd), .vdd(vdd), .A(_16847_), .B(_16842_), .C(_16848_), .Y(_16852_) );
	AND2X2 AND2X2_416 ( .gnd(gnd), .vdd(vdd), .A(_16600_), .B(_16583_), .Y(_16853_) );
	NAND3X1 NAND3X1_3476 ( .gnd(gnd), .vdd(vdd), .A(_16835_), .B(_16830_), .C(_16853_), .Y(_16855_) );
	NAND3X1 NAND3X1_3477 ( .gnd(gnd), .vdd(vdd), .A(_16852_), .B(_16855_), .C(_16851_), .Y(_16856_) );
	NAND3X1 NAND3X1_3478 ( .gnd(gnd), .vdd(vdd), .A(_16662_), .B(_16850_), .C(_16856_), .Y(_16857_) );
	INVX1 INVX1_2130 ( .gnd(gnd), .vdd(vdd), .A(_16597_), .Y(_16858_) );
	AOI21X1 AOI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_16608_), .B(_16604_), .C(_16858_), .Y(_16859_) );
	AOI21X1 AOI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_16855_), .B(_16852_), .C(_16851_), .Y(_16860_) );
	NOR3X1 NOR3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_16723_), .B(_16836_), .C(_16849_), .Y(_16861_) );
	OAI21X1 OAI21X1_3532 ( .gnd(gnd), .vdd(vdd), .A(_16861_), .B(_16860_), .C(_16859_), .Y(_16862_) );
	NAND3X1 NAND3X1_3479 ( .gnd(gnd), .vdd(vdd), .A(_16660_), .B(_16857_), .C(_16862_), .Y(_16863_) );
	OAI21X1 OAI21X1_3533 ( .gnd(gnd), .vdd(vdd), .A(_16861_), .B(_16860_), .C(_16662_), .Y(_16864_) );
	NAND3X1 NAND3X1_3480 ( .gnd(gnd), .vdd(vdd), .A(_16850_), .B(_16856_), .C(_16859_), .Y(_16866_) );
	NAND3X1 NAND3X1_3481 ( .gnd(gnd), .vdd(vdd), .A(_16659_), .B(_16866_), .C(_16864_), .Y(_16867_) );
	NAND3X1 NAND3X1_3482 ( .gnd(gnd), .vdd(vdd), .A(_16658_), .B(_16863_), .C(_16867_), .Y(_16868_) );
	AOI21X1 AOI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_16631_), .B(_16378_), .C(_16619_), .Y(_16869_) );
	NAND3X1 NAND3X1_3483 ( .gnd(gnd), .vdd(vdd), .A(_16659_), .B(_16857_), .C(_16862_), .Y(_16870_) );
	NAND3X1 NAND3X1_3484 ( .gnd(gnd), .vdd(vdd), .A(_16660_), .B(_16866_), .C(_16864_), .Y(_16871_) );
	NAND3X1 NAND3X1_3485 ( .gnd(gnd), .vdd(vdd), .A(_16869_), .B(_16870_), .C(_16871_), .Y(_16872_) );
	NAND2X1 NAND2X1_3360 ( .gnd(gnd), .vdd(vdd), .A(_16868_), .B(_16872_), .Y(_16873_) );
	NAND3X1 NAND3X1_3486 ( .gnd(gnd), .vdd(vdd), .A(_16628_), .B(_16631_), .C(_16630_), .Y(_16874_) );
	NAND2X1 NAND2X1_3361 ( .gnd(gnd), .vdd(vdd), .A(_16623_), .B(_16874_), .Y(_16875_) );
	AOI21X1 AOI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_16875_), .B(_16377_), .C(_16400_), .Y(_16877_) );
	NAND3X1 NAND3X1_3487 ( .gnd(gnd), .vdd(vdd), .A(_16378_), .B(_16631_), .C(_16630_), .Y(_16878_) );
	OAI21X1 OAI21X1_3534 ( .gnd(gnd), .vdd(vdd), .A(_16619_), .B(_16622_), .C(_16628_), .Y(_16879_) );
	NAND2X1 NAND2X1_3362 ( .gnd(gnd), .vdd(vdd), .A(_16879_), .B(_16878_), .Y(_16880_) );
	NOR3X1 NOR3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_16627_), .B(_16399_), .C(_16880_), .Y(_16881_) );
	OAI21X1 OAI21X1_3535 ( .gnd(gnd), .vdd(vdd), .A(_16877_), .B(_16881_), .C(_16873_), .Y(_16882_) );
	AND2X2 AND2X2_417 ( .gnd(gnd), .vdd(vdd), .A(_16872_), .B(_16868_), .Y(_16883_) );
	OAI21X1 OAI21X1_3536 ( .gnd(gnd), .vdd(vdd), .A(_16627_), .B(_16880_), .C(_16399_), .Y(_16884_) );
	NAND3X1 NAND3X1_3488 ( .gnd(gnd), .vdd(vdd), .A(_16377_), .B(_16400_), .C(_16875_), .Y(_16885_) );
	NAND3X1 NAND3X1_3489 ( .gnd(gnd), .vdd(vdd), .A(_16884_), .B(_16885_), .C(_16883_), .Y(_16886_) );
	NAND2X1 NAND2X1_3363 ( .gnd(gnd), .vdd(vdd), .A(_16882_), .B(_16886_), .Y(_16888_) );
	NAND3X1 NAND3X1_3490 ( .gnd(gnd), .vdd(vdd), .A(_16647_), .B(_16888_), .C(_16657_), .Y(_16889_) );
	OAI21X1 OAI21X1_3537 ( .gnd(gnd), .vdd(vdd), .A(_16877_), .B(_16881_), .C(_16883_), .Y(_16890_) );
	NAND3X1 NAND3X1_3491 ( .gnd(gnd), .vdd(vdd), .A(_16885_), .B(_16884_), .C(_16873_), .Y(_16891_) );
	NAND2X1 NAND2X1_3364 ( .gnd(gnd), .vdd(vdd), .A(_16891_), .B(_16890_), .Y(_16892_) );
	OAI21X1 OAI21X1_3538 ( .gnd(gnd), .vdd(vdd), .A(_16646_), .B(_16640_), .C(_16892_), .Y(_16893_) );
	NAND2X1 NAND2X1_3365 ( .gnd(gnd), .vdd(vdd), .A(_16889_), .B(_16893_), .Y(mulOut_31_) );
	NAND2X1 NAND2X1_3366 ( .gnd(gnd), .vdd(vdd), .A(_16722_), .B(_16799_), .Y(_16894_) );
	XNOR2X1 XNOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_16894_), .B(_15616_), .Y(mulOut_9_) );
	INVX1 INVX1_2131 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .Y(_17329_) );
	OAI21X1 OAI21X1_3539 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_1_), .B(pipelineStateController_pipelineState_0_), .C(_17329_), .Y(_17328__0_) );
	NAND2X1 NAND2X1_3367 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_0_), .B(_17329_), .Y(_17330_) );
	NOR2X1 NOR2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_1_), .B(_17330_), .Y(_17328__1_) );
	NAND2X1 NAND2X1_3368 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_1_), .B(_17329_), .Y(_17331_) );
	NOR2X1 NOR2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_0_), .B(_17331_), .Y(_17328__2_) );
	INVX1 INVX1_2132 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_1_), .Y(_17332_) );
	NOR2X1 NOR2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_17332_), .B(_17330_), .Y(_17328__3_) );
	OAI21X1 OAI21X1_3540 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_0_), .B(_427_), .C(_17329_), .Y(_17333_) );
	AOI21X1 AOI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_0_), .B(_427_), .C(_17333_), .Y(_17327__0_) );
	NAND2X1 NAND2X1_3369 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_0_), .B(_427_), .Y(_17334_) );
	NAND2X1 NAND2X1_3370 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_1_), .B(_17334_), .Y(_17335_) );
	NAND3X1 NAND3X1_3492 ( .gnd(gnd), .vdd(vdd), .A(pipelineStateController_pipelineState_0_), .B(_427_), .C(_17332_), .Y(_17336_) );
	AOI21X1 AOI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_17335_), .B(_17336_), .C(reset_bF_buf1), .Y(_17327__1_) );
	NOR2X1 NOR2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(executeState), .B(aOperand_we), .Y(_17337_) );
	OAI21X1 OAI21X1_3541 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(start), .C(aLoc_we), .Y(_17338_) );
	AOI21X1 AOI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_17338_), .B(_17337_), .C(reset_bF_buf0), .Y(_17326_) );
	DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17326_), .Q(_427_) );
	DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17327__0_), .Q(pipelineStateController_pipelineState_0_) );
	DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17327__1_), .Q(pipelineStateController_pipelineState_1_) );
	INVX1 INVX1_2133 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_2_), .Y(_17370_) );
	NOR3X1 NOR3X1_198 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(aLoc_frameOut_3_), .C(_17370_), .Y(_17371_) );
	INVX1 INVX1_2134 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .Y(_17372_) );
	NOR2X1 NOR2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_0_), .B(_17372_), .Y(_17373_) );
	NAND3X1 NAND3X1_3493 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_0_), .B(_17373__bF_buf5), .C(_17371__bF_buf7), .Y(_17374_) );
	NAND2X1 NAND2X1_3371 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .B(aLoc_frameOut_0_), .Y(_17375_) );
	INVX8 INVX8_72 ( .gnd(gnd), .vdd(vdd), .A(_17375_), .Y(_17376_) );
	NAND3X1 NAND3X1_3494 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_0_), .B(_17376__bF_buf5), .C(_17371__bF_buf6), .Y(_17377_) );
	NAND2X1 NAND2X1_3372 ( .gnd(gnd), .vdd(vdd), .A(_17374_), .B(_17377_), .Y(_17378_) );
	INVX1 INVX1_2135 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_0_), .Y(_17379_) );
	INVX1 INVX1_2136 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_0_), .Y(_17380_) );
	INVX4 INVX4_24 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .Y(_17381_) );
	NOR2X1 NOR2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_3_), .B(aLoc_frameOut_2_), .Y(_17382_) );
	NAND3X1 NAND3X1_3495 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17382_), .C(_17373__bF_buf4), .Y(_17383_) );
	NAND3X1 NAND3X1_3496 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17382_), .C(_17376__bF_buf4), .Y(_17384_) );
	OAI22X1 OAI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(_17379_), .B(_17384__bF_buf4), .C(_17380_), .D(_17383__bF_buf4), .Y(_17385_) );
	NOR2X1 NOR2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_17378_), .B(_17385_), .Y(_17386_) );
	INVX1 INVX1_2137 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_0_), .Y(_17387_) );
	INVX1 INVX1_2138 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_0_), .Y(_17388_) );
	INVX1 INVX1_2139 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_0_), .Y(_17389_) );
	NOR2X1 NOR2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .B(_17389_), .Y(_17390_) );
	INVX1 INVX1_2140 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_3_), .Y(_17391_) );
	NOR2X1 NOR2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_2_), .B(_17391_), .Y(_17392_) );
	NAND3X1 NAND3X1_3497 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17390_), .C(_17392__bF_buf7), .Y(_17393_) );
	NAND3X1 NAND3X1_3498 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17376__bF_buf3), .C(_17392__bF_buf6), .Y(_17394_) );
	OAI22X1 OAI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(_17387_), .B(_17394__bF_buf4), .C(_17388_), .D(_17393__bF_buf4), .Y(_17395_) );
	INVX1 INVX1_2141 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_0_), .Y(_17396_) );
	INVX1 INVX1_2142 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_0_), .Y(_17397_) );
	NAND2X1 NAND2X1_3373 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_3_), .B(aLoc_frameOut_2_), .Y(_17398_) );
	INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(_17398_), .Y(_17399_) );
	NAND3X1 NAND3X1_3499 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17399_), .C(_17390_), .Y(_17400_) );
	NAND3X1 NAND3X1_3500 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17399_), .C(_17373__bF_buf3), .Y(_17401_) );
	OAI22X1 OAI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(_17396_), .B(_17401__bF_buf4), .C(_17397_), .D(_17400__bF_buf4), .Y(_17402_) );
	NOR2X1 NOR2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_17402_), .B(_17395_), .Y(_17403_) );
	NAND2X1 NAND2X1_3374 ( .gnd(gnd), .vdd(vdd), .A(_17386_), .B(_17403_), .Y(_17404_) );
	INVX1 INVX1_2143 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_0_), .Y(_17405_) );
	INVX1 INVX1_2144 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_0_), .Y(_17406_) );
	NAND3X1 NAND3X1_3501 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(_17382_), .C(_17373__bF_buf2), .Y(_17407_) );
	NAND3X1 NAND3X1_3502 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(_17382_), .C(_17376__bF_buf2), .Y(_17408_) );
	OAI22X1 OAI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_17406_), .B(_17408__bF_buf4), .C(_17405_), .D(_17407__bF_buf4), .Y(_17409_) );
	INVX1 INVX1_2145 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_0_), .Y(_17410_) );
	NOR2X1 NOR2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_3_), .B(_17370_), .Y(_17411_) );
	NAND3X1 NAND3X1_3503 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(_17390_), .C(_17411__bF_buf5), .Y(_17412_) );
	NOR3X1 NOR3X1_199 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .B(aLoc_frameOut_0_), .C(_17381_), .Y(_17413_) );
	NAND3X1 NAND3X1_3504 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_0_), .B(_17411__bF_buf4), .C(_17413__bF_buf7), .Y(_17414_) );
	OAI21X1 OAI21X1_3542 ( .gnd(gnd), .vdd(vdd), .A(_17410_), .B(_17412__bF_buf4), .C(_17414_), .Y(_17415_) );
	NOR2X1 NOR2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_17409_), .B(_17415_), .Y(_17416_) );
	INVX1 INVX1_2146 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_0_), .Y(_17417_) );
	NAND3X1 NAND3X1_3505 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(_17399_), .C(_17373__bF_buf1), .Y(_17418_) );
	NOR2X1 NOR2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_17398_), .B(_17375_), .Y(_17419_) );
	NAND3X1 NAND3X1_3506 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(registers_r31_0_), .C(_17419__bF_buf4), .Y(_17420_) );
	OAI21X1 OAI21X1_3543 ( .gnd(gnd), .vdd(vdd), .A(_17417_), .B(_17418__bF_buf4), .C(_17420_), .Y(_17421_) );
	INVX1 INVX1_2147 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_0_), .Y(_17422_) );
	NAND3X1 NAND3X1_3507 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(_17390_), .C(_17392__bF_buf5), .Y(_17423_) );
	NAND3X1 NAND3X1_3508 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_0_), .B(_17392__bF_buf4), .C(_17413__bF_buf6), .Y(_17424_) );
	OAI21X1 OAI21X1_3544 ( .gnd(gnd), .vdd(vdd), .A(_17422_), .B(_17423__bF_buf4), .C(_17424_), .Y(_17425_) );
	NOR2X1 NOR2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_17421_), .B(_17425_), .Y(_17426_) );
	NAND2X1 NAND2X1_3375 ( .gnd(gnd), .vdd(vdd), .A(_17426_), .B(_17416_), .Y(_17427_) );
	NOR2X1 NOR2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_17427_), .B(_17404_), .Y(_17428_) );
	NAND2X1 NAND2X1_3376 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_0_), .B(_17372_), .Y(_17429_) );
	INVX1 INVX1_2148 ( .gnd(gnd), .vdd(vdd), .A(_17382_), .Y(_17430_) );
	NOR3X1 NOR3X1_200 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .B(_17429_), .C(_17430_), .Y(_17431_) );
	NOR3X1 NOR3X1_201 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(aLoc_frameOut_1_), .C(aLoc_frameOut_0_), .Y(_17432_) );
	AND2X2 AND2X2_418 ( .gnd(gnd), .vdd(vdd), .A(_17432__bF_buf4), .B(_17399_), .Y(_17433_) );
	AOI22X1 AOI22X1_378 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_0_), .C(registers_r1_0_), .D(_17431__bF_buf4), .Y(_17434_) );
	AND2X2 AND2X2_419 ( .gnd(gnd), .vdd(vdd), .A(_17411__bF_buf3), .B(_17432__bF_buf3), .Y(_17435_) );
	AND2X2 AND2X2_420 ( .gnd(gnd), .vdd(vdd), .A(_17371__bF_buf5), .B(_17390_), .Y(_17436_) );
	AOI22X1 AOI22X1_379 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_0_), .C(registers_r5_0_), .D(_17436__bF_buf4), .Y(_17437_) );
	NAND2X1 NAND2X1_3377 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .B(_17389_), .Y(_17438_) );
	NAND2X1 NAND2X1_3378 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_3_), .B(_17370_), .Y(_17439_) );
	NOR3X1 NOR3X1_202 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(_17438_), .C(_17439_), .Y(_17440_) );
	INVX1 INVX1_2149 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_0_), .Y(_17441_) );
	NAND3X1 NAND3X1_3509 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_0_), .B(_17432__bF_buf2), .C(_17392__bF_buf3), .Y(_17442_) );
	NAND3X1 NAND3X1_3510 ( .gnd(gnd), .vdd(vdd), .A(_17381_), .B(_17399_), .C(_17376__bF_buf1), .Y(_17443_) );
	OAI21X1 OAI21X1_3545 ( .gnd(gnd), .vdd(vdd), .A(_17441_), .B(_17443__bF_buf4), .C(_17442_), .Y(_17444_) );
	AOI21X1 AOI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_0_), .B(_17440__bF_buf4), .C(_17444_), .Y(_17445_) );
	NAND3X1 NAND3X1_3511 ( .gnd(gnd), .vdd(vdd), .A(_17434_), .B(_17437_), .C(_17445_), .Y(_17446_) );
	INVX1 INVX1_2150 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_0_), .Y(_17447_) );
	INVX1 INVX1_2151 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_0_), .Y(_17448_) );
	NAND3X1 NAND3X1_3512 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(_17411__bF_buf2), .C(_17373__bF_buf0), .Y(_17449_) );
	NAND3X1 NAND3X1_3513 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(_17376__bF_buf0), .C(_17411__bF_buf1), .Y(_17450_) );
	OAI22X1 OAI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(_17448_), .B(_17450__bF_buf4), .C(_17447_), .D(_17449__bF_buf4), .Y(_17451_) );
	INVX1 INVX1_2152 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_0_), .Y(_17452_) );
	INVX1 INVX1_2153 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_0_), .Y(_17453_) );
	NAND3X1 NAND3X1_3514 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(_17382_), .C(_17390_), .Y(_17454_) );
	NOR2X1 NOR2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_1_), .B(aLoc_frameOut_0_), .Y(_17455_) );
	NAND3X1 NAND3X1_3515 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(_17382_), .C(_17455_), .Y(_17456_) );
	OAI22X1 OAI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(_17452_), .B(_17456__bF_buf4), .C(_17453_), .D(_17454__bF_buf4), .Y(_17457_) );
	NOR2X1 NOR2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_17457_), .B(_17451_), .Y(_17458_) );
	INVX1 INVX1_2154 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_0_), .Y(_17459_) );
	INVX1 INVX1_2155 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_0_), .Y(_17460_) );
	NAND3X1 NAND3X1_3516 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .B(_17455_), .C(_17399_), .Y(_17461_) );
	NAND3X1 NAND3X1_3517 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(_17399_), .C(_17390_), .Y(_17462_) );
	OAI22X1 OAI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(_17459_), .B(_17461__bF_buf4), .C(_17460_), .D(_17462__bF_buf4), .Y(_17463_) );
	INVX1 INVX1_2156 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_0_), .Y(_17464_) );
	INVX1 INVX1_2157 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_0_), .Y(_17465_) );
	NAND3X1 NAND3X1_3518 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(_17373__bF_buf5), .C(_17392__bF_buf2), .Y(_17466_) );
	NAND3X1 NAND3X1_3519 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(_17376__bF_buf5), .C(_17392__bF_buf1), .Y(_17467_) );
	OAI22X1 OAI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(_17465_), .B(_17467__bF_buf4), .C(_17464_), .D(_17466__bF_buf4), .Y(_17468_) );
	NOR2X1 NOR2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_17463_), .B(_17468_), .Y(_17469_) );
	NAND2X1 NAND2X1_3379 ( .gnd(gnd), .vdd(vdd), .A(_17458_), .B(_17469_), .Y(_17470_) );
	NOR2X1 NOR2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_17446_), .B(_17470_), .Y(_17471_) );
	NAND2X1 NAND2X1_3380 ( .gnd(gnd), .vdd(vdd), .A(_17471_), .B(_17428_), .Y(_428__0_) );
	NAND3X1 NAND3X1_3520 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_1_), .B(_17373__bF_buf4), .C(_17371__bF_buf4), .Y(_17472_) );
	NAND3X1 NAND3X1_3521 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_1_), .B(_17376__bF_buf4), .C(_17371__bF_buf3), .Y(_17473_) );
	NAND2X1 NAND2X1_3381 ( .gnd(gnd), .vdd(vdd), .A(_17472_), .B(_17473_), .Y(_17474_) );
	INVX1 INVX1_2158 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_1_), .Y(_17475_) );
	INVX1 INVX1_2159 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_1_), .Y(_17476_) );
	OAI22X1 OAI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(_17475_), .B(_17384__bF_buf3), .C(_17476_), .D(_17383__bF_buf3), .Y(_17477_) );
	NOR2X1 NOR2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_17474_), .B(_17477_), .Y(_17478_) );
	INVX1 INVX1_2160 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_1_), .Y(_17479_) );
	INVX1 INVX1_2161 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_1_), .Y(_17480_) );
	OAI22X1 OAI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(_17479_), .B(_17394__bF_buf3), .C(_17480_), .D(_17393__bF_buf3), .Y(_17481_) );
	INVX1 INVX1_2162 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_1_), .Y(_17482_) );
	INVX1 INVX1_2163 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_1_), .Y(_17483_) );
	OAI22X1 OAI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(_17482_), .B(_17401__bF_buf3), .C(_17483_), .D(_17400__bF_buf3), .Y(_17484_) );
	NOR2X1 NOR2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_17484_), .B(_17481_), .Y(_17485_) );
	NAND2X1 NAND2X1_3382 ( .gnd(gnd), .vdd(vdd), .A(_17478_), .B(_17485_), .Y(_17486_) );
	INVX1 INVX1_2164 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_1_), .Y(_17487_) );
	INVX1 INVX1_2165 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_1_), .Y(_17488_) );
	OAI22X1 OAI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(_17488_), .B(_17408__bF_buf3), .C(_17487_), .D(_17407__bF_buf3), .Y(_17489_) );
	INVX1 INVX1_2166 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_1_), .Y(_17490_) );
	NAND3X1 NAND3X1_3522 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_1_), .B(_17411__bF_buf0), .C(_17413__bF_buf5), .Y(_17491_) );
	OAI21X1 OAI21X1_3546 ( .gnd(gnd), .vdd(vdd), .A(_17490_), .B(_17412__bF_buf3), .C(_17491_), .Y(_17492_) );
	NOR2X1 NOR2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_17489_), .B(_17492_), .Y(_17493_) );
	INVX1 INVX1_2167 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_1_), .Y(_17494_) );
	NAND3X1 NAND3X1_3523 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(registers_r31_1_), .C(_17419__bF_buf3), .Y(_17495_) );
	OAI21X1 OAI21X1_3547 ( .gnd(gnd), .vdd(vdd), .A(_17494_), .B(_17418__bF_buf3), .C(_17495_), .Y(_17496_) );
	INVX1 INVX1_2168 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_1_), .Y(_17497_) );
	NAND3X1 NAND3X1_3524 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_1_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_17498_) );
	OAI21X1 OAI21X1_3548 ( .gnd(gnd), .vdd(vdd), .A(_17497_), .B(_17423__bF_buf3), .C(_17498_), .Y(_17499_) );
	NOR2X1 NOR2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_17496_), .B(_17499_), .Y(_17500_) );
	NAND2X1 NAND2X1_3383 ( .gnd(gnd), .vdd(vdd), .A(_17500_), .B(_17493_), .Y(_17501_) );
	NOR2X1 NOR2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_17501_), .B(_17486_), .Y(_17502_) );
	AOI22X1 AOI22X1_380 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_1_), .C(registers_r1_1_), .D(_17431__bF_buf3), .Y(_17503_) );
	AOI22X1 AOI22X1_381 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_1_), .C(registers_r5_1_), .D(_17436__bF_buf3), .Y(_17504_) );
	INVX1 INVX1_2169 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_1_), .Y(_17505_) );
	NAND3X1 NAND3X1_3525 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_1_), .B(_17432__bF_buf1), .C(_17392__bF_buf7), .Y(_17506_) );
	OAI21X1 OAI21X1_3549 ( .gnd(gnd), .vdd(vdd), .A(_17505_), .B(_17443__bF_buf3), .C(_17506_), .Y(_17507_) );
	AOI21X1 AOI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_1_), .B(_17440__bF_buf3), .C(_17507_), .Y(_17508_) );
	NAND3X1 NAND3X1_3526 ( .gnd(gnd), .vdd(vdd), .A(_17503_), .B(_17504_), .C(_17508_), .Y(_17509_) );
	INVX1 INVX1_2170 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_1_), .Y(_17510_) );
	INVX1 INVX1_2171 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_1_), .Y(_17511_) );
	OAI22X1 OAI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(_17511_), .B(_17450__bF_buf3), .C(_17510_), .D(_17449__bF_buf3), .Y(_17512_) );
	INVX1 INVX1_2172 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_1_), .Y(_17513_) );
	INVX1 INVX1_2173 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_1_), .Y(_17514_) );
	OAI22X1 OAI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(_17513_), .B(_17456__bF_buf3), .C(_17514_), .D(_17454__bF_buf3), .Y(_17515_) );
	NOR2X1 NOR2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_17515_), .B(_17512_), .Y(_17516_) );
	INVX1 INVX1_2174 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_1_), .Y(_17517_) );
	INVX1 INVX1_2175 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_1_), .Y(_17518_) );
	OAI22X1 OAI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(_17517_), .B(_17461__bF_buf3), .C(_17518_), .D(_17462__bF_buf3), .Y(_17519_) );
	INVX1 INVX1_2176 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_1_), .Y(_17520_) );
	INVX1 INVX1_2177 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_1_), .Y(_17521_) );
	OAI22X1 OAI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(_17521_), .B(_17467__bF_buf3), .C(_17520_), .D(_17466__bF_buf3), .Y(_17522_) );
	NOR2X1 NOR2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_17519_), .B(_17522_), .Y(_17523_) );
	NAND2X1 NAND2X1_3384 ( .gnd(gnd), .vdd(vdd), .A(_17516_), .B(_17523_), .Y(_17524_) );
	NOR2X1 NOR2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_17509_), .B(_17524_), .Y(_17525_) );
	NAND2X1 NAND2X1_3385 ( .gnd(gnd), .vdd(vdd), .A(_17525_), .B(_17502_), .Y(_428__1_) );
	NAND3X1 NAND3X1_3527 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_2_), .B(_17373__bF_buf3), .C(_17371__bF_buf2), .Y(_17526_) );
	NAND3X1 NAND3X1_3528 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_2_), .B(_17376__bF_buf3), .C(_17371__bF_buf1), .Y(_17527_) );
	NAND2X1 NAND2X1_3386 ( .gnd(gnd), .vdd(vdd), .A(_17526_), .B(_17527_), .Y(_17528_) );
	INVX1 INVX1_2178 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_2_), .Y(_17529_) );
	INVX1 INVX1_2179 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_2_), .Y(_17530_) );
	OAI22X1 OAI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(_17529_), .B(_17384__bF_buf2), .C(_17530_), .D(_17383__bF_buf2), .Y(_17531_) );
	NOR2X1 NOR2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_17528_), .B(_17531_), .Y(_17532_) );
	INVX1 INVX1_2180 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_2_), .Y(_17533_) );
	INVX1 INVX1_2181 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_2_), .Y(_17534_) );
	OAI22X1 OAI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(_17533_), .B(_17394__bF_buf2), .C(_17534_), .D(_17393__bF_buf2), .Y(_17535_) );
	INVX1 INVX1_2182 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_2_), .Y(_17536_) );
	INVX1 INVX1_2183 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_2_), .Y(_17537_) );
	OAI22X1 OAI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(_17536_), .B(_17401__bF_buf2), .C(_17537_), .D(_17400__bF_buf2), .Y(_17538_) );
	NOR2X1 NOR2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_17538_), .B(_17535_), .Y(_17539_) );
	NAND2X1 NAND2X1_3387 ( .gnd(gnd), .vdd(vdd), .A(_17532_), .B(_17539_), .Y(_17540_) );
	INVX1 INVX1_2184 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_2_), .Y(_17541_) );
	INVX1 INVX1_2185 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_2_), .Y(_17542_) );
	OAI22X1 OAI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(_17542_), .B(_17408__bF_buf2), .C(_17541_), .D(_17407__bF_buf2), .Y(_17543_) );
	INVX1 INVX1_2186 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_2_), .Y(_17544_) );
	NAND3X1 NAND3X1_3529 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_2_), .B(_17411__bF_buf5), .C(_17413__bF_buf3), .Y(_17545_) );
	OAI21X1 OAI21X1_3550 ( .gnd(gnd), .vdd(vdd), .A(_17544_), .B(_17412__bF_buf2), .C(_17545_), .Y(_17546_) );
	NOR2X1 NOR2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_17543_), .B(_17546_), .Y(_17547_) );
	INVX1 INVX1_2187 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_2_), .Y(_17548_) );
	NAND3X1 NAND3X1_3530 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(registers_r31_2_), .C(_17419__bF_buf2), .Y(_17549_) );
	OAI21X1 OAI21X1_3551 ( .gnd(gnd), .vdd(vdd), .A(_17548_), .B(_17418__bF_buf2), .C(_17549_), .Y(_17550_) );
	INVX1 INVX1_2188 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_2_), .Y(_17551_) );
	NAND3X1 NAND3X1_3531 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_2_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_17552_) );
	OAI21X1 OAI21X1_3552 ( .gnd(gnd), .vdd(vdd), .A(_17551_), .B(_17423__bF_buf2), .C(_17552_), .Y(_17553_) );
	NOR2X1 NOR2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_17550_), .B(_17553_), .Y(_17554_) );
	NAND2X1 NAND2X1_3388 ( .gnd(gnd), .vdd(vdd), .A(_17554_), .B(_17547_), .Y(_17555_) );
	NOR2X1 NOR2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_17555_), .B(_17540_), .Y(_17556_) );
	AOI22X1 AOI22X1_382 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf2), .B(registers_a2_2_), .C(registers_r1_2_), .D(_17431__bF_buf2), .Y(_17557_) );
	AOI22X1 AOI22X1_383 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf2), .B(registers_r4_2_), .C(registers_r5_2_), .D(_17436__bF_buf2), .Y(_17558_) );
	INVX1 INVX1_2189 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_2_), .Y(_17559_) );
	NAND3X1 NAND3X1_3532 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_2_), .B(_17432__bF_buf0), .C(_17392__bF_buf5), .Y(_17560_) );
	OAI21X1 OAI21X1_3553 ( .gnd(gnd), .vdd(vdd), .A(_17559_), .B(_17443__bF_buf2), .C(_17560_), .Y(_17561_) );
	AOI21X1 AOI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_2_), .B(_17440__bF_buf2), .C(_17561_), .Y(_17562_) );
	NAND3X1 NAND3X1_3533 ( .gnd(gnd), .vdd(vdd), .A(_17557_), .B(_17558_), .C(_17562_), .Y(_17563_) );
	INVX1 INVX1_2190 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_2_), .Y(_17564_) );
	INVX1 INVX1_2191 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_2_), .Y(_17565_) );
	OAI22X1 OAI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(_17565_), .B(_17450__bF_buf2), .C(_17564_), .D(_17449__bF_buf2), .Y(_17566_) );
	INVX1 INVX1_2192 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_2_), .Y(_17567_) );
	INVX1 INVX1_2193 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_2_), .Y(_17568_) );
	OAI22X1 OAI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(_17567_), .B(_17456__bF_buf2), .C(_17568_), .D(_17454__bF_buf2), .Y(_17569_) );
	NOR2X1 NOR2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_17569_), .B(_17566_), .Y(_17570_) );
	INVX1 INVX1_2194 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_2_), .Y(_17571_) );
	INVX1 INVX1_2195 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_2_), .Y(_17572_) );
	OAI22X1 OAI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(_17571_), .B(_17461__bF_buf2), .C(_17572_), .D(_17462__bF_buf2), .Y(_17573_) );
	INVX1 INVX1_2196 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_2_), .Y(_17574_) );
	INVX1 INVX1_2197 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_2_), .Y(_17575_) );
	OAI22X1 OAI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(_17575_), .B(_17467__bF_buf2), .C(_17574_), .D(_17466__bF_buf2), .Y(_17576_) );
	NOR2X1 NOR2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_17573_), .B(_17576_), .Y(_17577_) );
	NAND2X1 NAND2X1_3389 ( .gnd(gnd), .vdd(vdd), .A(_17570_), .B(_17577_), .Y(_17578_) );
	NOR2X1 NOR2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_17563_), .B(_17578_), .Y(_17579_) );
	NAND2X1 NAND2X1_3390 ( .gnd(gnd), .vdd(vdd), .A(_17579_), .B(_17556_), .Y(_428__2_) );
	NAND3X1 NAND3X1_3534 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_3_), .B(_17373__bF_buf2), .C(_17371__bF_buf0), .Y(_17580_) );
	NAND3X1 NAND3X1_3535 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_3_), .B(_17376__bF_buf2), .C(_17371__bF_buf7), .Y(_17581_) );
	NAND2X1 NAND2X1_3391 ( .gnd(gnd), .vdd(vdd), .A(_17580_), .B(_17581_), .Y(_17582_) );
	INVX1 INVX1_2198 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_3_), .Y(_17583_) );
	INVX1 INVX1_2199 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_3_), .Y(_17584_) );
	OAI22X1 OAI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(_17583_), .B(_17384__bF_buf1), .C(_17584_), .D(_17383__bF_buf1), .Y(_17585_) );
	NOR2X1 NOR2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_17582_), .B(_17585_), .Y(_17586_) );
	INVX1 INVX1_2200 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_3_), .Y(_17587_) );
	INVX1 INVX1_2201 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_3_), .Y(_17588_) );
	OAI22X1 OAI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(_17587_), .B(_17394__bF_buf1), .C(_17588_), .D(_17393__bF_buf1), .Y(_17589_) );
	INVX1 INVX1_2202 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_3_), .Y(_17590_) );
	INVX1 INVX1_2203 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_3_), .Y(_17591_) );
	OAI22X1 OAI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(_17590_), .B(_17401__bF_buf1), .C(_17591_), .D(_17400__bF_buf1), .Y(_17592_) );
	NOR2X1 NOR2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_17592_), .B(_17589_), .Y(_17593_) );
	NAND2X1 NAND2X1_3392 ( .gnd(gnd), .vdd(vdd), .A(_17586_), .B(_17593_), .Y(_17594_) );
	INVX1 INVX1_2204 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_3_), .Y(_17595_) );
	INVX1 INVX1_2205 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_3_), .Y(_17596_) );
	OAI22X1 OAI22X1_179 ( .gnd(gnd), .vdd(vdd), .A(_17596_), .B(_17408__bF_buf1), .C(_17595_), .D(_17407__bF_buf1), .Y(_17597_) );
	INVX1 INVX1_2206 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_3_), .Y(_17598_) );
	NAND3X1 NAND3X1_3536 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_3_), .B(_17411__bF_buf4), .C(_17413__bF_buf1), .Y(_17599_) );
	OAI21X1 OAI21X1_3554 ( .gnd(gnd), .vdd(vdd), .A(_17598_), .B(_17412__bF_buf1), .C(_17599_), .Y(_17600_) );
	NOR2X1 NOR2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_17597_), .B(_17600_), .Y(_17601_) );
	INVX1 INVX1_2207 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_3_), .Y(_17602_) );
	NAND3X1 NAND3X1_3537 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(registers_r31_3_), .C(_17419__bF_buf1), .Y(_17603_) );
	OAI21X1 OAI21X1_3555 ( .gnd(gnd), .vdd(vdd), .A(_17602_), .B(_17418__bF_buf1), .C(_17603_), .Y(_17604_) );
	INVX1 INVX1_2208 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_3_), .Y(_17605_) );
	NAND3X1 NAND3X1_3538 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_3_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_17606_) );
	OAI21X1 OAI21X1_3556 ( .gnd(gnd), .vdd(vdd), .A(_17605_), .B(_17423__bF_buf1), .C(_17606_), .Y(_17607_) );
	NOR2X1 NOR2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_17604_), .B(_17607_), .Y(_17608_) );
	NAND2X1 NAND2X1_3393 ( .gnd(gnd), .vdd(vdd), .A(_17608_), .B(_17601_), .Y(_17609_) );
	NOR2X1 NOR2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_17609_), .B(_17594_), .Y(_17610_) );
	AOI22X1 AOI22X1_384 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf1), .B(registers_a2_3_), .C(registers_r1_3_), .D(_17431__bF_buf1), .Y(_17611_) );
	AOI22X1 AOI22X1_385 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf1), .B(registers_r4_3_), .C(registers_r5_3_), .D(_17436__bF_buf1), .Y(_17612_) );
	INVX1 INVX1_2209 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_3_), .Y(_17613_) );
	NAND3X1 NAND3X1_3539 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_3_), .B(_17432__bF_buf4), .C(_17392__bF_buf3), .Y(_17614_) );
	OAI21X1 OAI21X1_3557 ( .gnd(gnd), .vdd(vdd), .A(_17613_), .B(_17443__bF_buf1), .C(_17614_), .Y(_17615_) );
	AOI21X1 AOI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_3_), .B(_17440__bF_buf1), .C(_17615_), .Y(_17616_) );
	NAND3X1 NAND3X1_3540 ( .gnd(gnd), .vdd(vdd), .A(_17611_), .B(_17612_), .C(_17616_), .Y(_17617_) );
	INVX1 INVX1_2210 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_3_), .Y(_17618_) );
	INVX1 INVX1_2211 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_3_), .Y(_17619_) );
	OAI22X1 OAI22X1_180 ( .gnd(gnd), .vdd(vdd), .A(_17619_), .B(_17450__bF_buf1), .C(_17618_), .D(_17449__bF_buf1), .Y(_17620_) );
	INVX1 INVX1_2212 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_3_), .Y(_17621_) );
	INVX1 INVX1_2213 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_3_), .Y(_17622_) );
	OAI22X1 OAI22X1_181 ( .gnd(gnd), .vdd(vdd), .A(_17621_), .B(_17456__bF_buf1), .C(_17622_), .D(_17454__bF_buf1), .Y(_17623_) );
	NOR2X1 NOR2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_17623_), .B(_17620_), .Y(_17624_) );
	INVX1 INVX1_2214 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_3_), .Y(_17625_) );
	INVX1 INVX1_2215 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_3_), .Y(_17626_) );
	OAI22X1 OAI22X1_182 ( .gnd(gnd), .vdd(vdd), .A(_17625_), .B(_17461__bF_buf1), .C(_17626_), .D(_17462__bF_buf1), .Y(_17627_) );
	INVX1 INVX1_2216 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_3_), .Y(_17628_) );
	INVX1 INVX1_2217 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_3_), .Y(_17629_) );
	OAI22X1 OAI22X1_183 ( .gnd(gnd), .vdd(vdd), .A(_17629_), .B(_17467__bF_buf1), .C(_17628_), .D(_17466__bF_buf1), .Y(_17630_) );
	NOR2X1 NOR2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_17627_), .B(_17630_), .Y(_17631_) );
	NAND2X1 NAND2X1_3394 ( .gnd(gnd), .vdd(vdd), .A(_17624_), .B(_17631_), .Y(_17632_) );
	NOR2X1 NOR2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_17617_), .B(_17632_), .Y(_17633_) );
	NAND2X1 NAND2X1_3395 ( .gnd(gnd), .vdd(vdd), .A(_17633_), .B(_17610_), .Y(_428__3_) );
	NAND3X1 NAND3X1_3541 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_4_), .B(_17373__bF_buf1), .C(_17371__bF_buf6), .Y(_17634_) );
	NAND3X1 NAND3X1_3542 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_4_), .B(_17376__bF_buf1), .C(_17371__bF_buf5), .Y(_17635_) );
	NAND2X1 NAND2X1_3396 ( .gnd(gnd), .vdd(vdd), .A(_17634_), .B(_17635_), .Y(_17636_) );
	INVX1 INVX1_2218 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_4_), .Y(_17637_) );
	INVX1 INVX1_2219 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_4_), .Y(_17638_) );
	OAI22X1 OAI22X1_184 ( .gnd(gnd), .vdd(vdd), .A(_17637_), .B(_17384__bF_buf0), .C(_17638_), .D(_17383__bF_buf0), .Y(_17639_) );
	NOR2X1 NOR2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_17636_), .B(_17639_), .Y(_17640_) );
	INVX1 INVX1_2220 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_4_), .Y(_17641_) );
	INVX1 INVX1_2221 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_4_), .Y(_17642_) );
	OAI22X1 OAI22X1_185 ( .gnd(gnd), .vdd(vdd), .A(_17641_), .B(_17394__bF_buf0), .C(_17642_), .D(_17393__bF_buf0), .Y(_17643_) );
	INVX1 INVX1_2222 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_4_), .Y(_17644_) );
	INVX1 INVX1_2223 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_4_), .Y(_17645_) );
	OAI22X1 OAI22X1_186 ( .gnd(gnd), .vdd(vdd), .A(_17644_), .B(_17401__bF_buf0), .C(_17645_), .D(_17400__bF_buf0), .Y(_17646_) );
	NOR2X1 NOR2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_17646_), .B(_17643_), .Y(_17647_) );
	NAND2X1 NAND2X1_3397 ( .gnd(gnd), .vdd(vdd), .A(_17640_), .B(_17647_), .Y(_17648_) );
	INVX1 INVX1_2224 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_4_), .Y(_17649_) );
	INVX1 INVX1_2225 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_4_), .Y(_17650_) );
	OAI22X1 OAI22X1_187 ( .gnd(gnd), .vdd(vdd), .A(_17650_), .B(_17408__bF_buf0), .C(_17649_), .D(_17407__bF_buf0), .Y(_17651_) );
	INVX1 INVX1_2226 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_4_), .Y(_17652_) );
	NAND3X1 NAND3X1_3543 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_4_), .B(_17411__bF_buf3), .C(_17413__bF_buf7), .Y(_17653_) );
	OAI21X1 OAI21X1_3558 ( .gnd(gnd), .vdd(vdd), .A(_17652_), .B(_17412__bF_buf0), .C(_17653_), .Y(_17654_) );
	NOR2X1 NOR2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_17651_), .B(_17654_), .Y(_17655_) );
	INVX1 INVX1_2227 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_4_), .Y(_17656_) );
	NAND3X1 NAND3X1_3544 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .B(registers_r31_4_), .C(_17419__bF_buf0), .Y(_17657_) );
	OAI21X1 OAI21X1_3559 ( .gnd(gnd), .vdd(vdd), .A(_17656_), .B(_17418__bF_buf0), .C(_17657_), .Y(_17658_) );
	INVX1 INVX1_2228 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_4_), .Y(_17659_) );
	NAND3X1 NAND3X1_3545 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_4_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_17660_) );
	OAI21X1 OAI21X1_3560 ( .gnd(gnd), .vdd(vdd), .A(_17659_), .B(_17423__bF_buf0), .C(_17660_), .Y(_17661_) );
	NOR2X1 NOR2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_17658_), .B(_17661_), .Y(_17662_) );
	NAND2X1 NAND2X1_3398 ( .gnd(gnd), .vdd(vdd), .A(_17662_), .B(_17655_), .Y(_17663_) );
	NOR2X1 NOR2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_17663_), .B(_17648_), .Y(_17664_) );
	AOI22X1 AOI22X1_386 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf0), .B(registers_a2_4_), .C(registers_r1_4_), .D(_17431__bF_buf0), .Y(_17665_) );
	AOI22X1 AOI22X1_387 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf0), .B(registers_r4_4_), .C(registers_r5_4_), .D(_17436__bF_buf0), .Y(_17666_) );
	INVX1 INVX1_2229 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_4_), .Y(_17667_) );
	NAND3X1 NAND3X1_3546 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_4_), .B(_17432__bF_buf3), .C(_17392__bF_buf1), .Y(_17668_) );
	OAI21X1 OAI21X1_3561 ( .gnd(gnd), .vdd(vdd), .A(_17667_), .B(_17443__bF_buf0), .C(_17668_), .Y(_17669_) );
	AOI21X1 AOI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_4_), .B(_17440__bF_buf0), .C(_17669_), .Y(_17670_) );
	NAND3X1 NAND3X1_3547 ( .gnd(gnd), .vdd(vdd), .A(_17665_), .B(_17666_), .C(_17670_), .Y(_17671_) );
	INVX1 INVX1_2230 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_4_), .Y(_17672_) );
	INVX1 INVX1_2231 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_4_), .Y(_17673_) );
	OAI22X1 OAI22X1_188 ( .gnd(gnd), .vdd(vdd), .A(_17673_), .B(_17450__bF_buf0), .C(_17672_), .D(_17449__bF_buf0), .Y(_17674_) );
	INVX1 INVX1_2232 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_4_), .Y(_17675_) );
	INVX1 INVX1_2233 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_4_), .Y(_17676_) );
	OAI22X1 OAI22X1_189 ( .gnd(gnd), .vdd(vdd), .A(_17675_), .B(_17456__bF_buf0), .C(_17676_), .D(_17454__bF_buf0), .Y(_17677_) );
	NOR2X1 NOR2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_17677_), .B(_17674_), .Y(_17678_) );
	INVX1 INVX1_2234 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_4_), .Y(_17679_) );
	INVX1 INVX1_2235 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_4_), .Y(_17680_) );
	OAI22X1 OAI22X1_190 ( .gnd(gnd), .vdd(vdd), .A(_17679_), .B(_17461__bF_buf0), .C(_17680_), .D(_17462__bF_buf0), .Y(_17681_) );
	INVX1 INVX1_2236 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_4_), .Y(_17682_) );
	INVX1 INVX1_2237 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_4_), .Y(_17683_) );
	OAI22X1 OAI22X1_191 ( .gnd(gnd), .vdd(vdd), .A(_17683_), .B(_17467__bF_buf0), .C(_17682_), .D(_17466__bF_buf0), .Y(_17684_) );
	NOR2X1 NOR2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_17681_), .B(_17684_), .Y(_17685_) );
	NAND2X1 NAND2X1_3399 ( .gnd(gnd), .vdd(vdd), .A(_17678_), .B(_17685_), .Y(_17686_) );
	NOR2X1 NOR2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_17671_), .B(_17686_), .Y(_17687_) );
	NAND2X1 NAND2X1_3400 ( .gnd(gnd), .vdd(vdd), .A(_17687_), .B(_17664_), .Y(_428__4_) );
	NAND3X1 NAND3X1_3548 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_5_), .B(_17373__bF_buf0), .C(_17371__bF_buf4), .Y(_17688_) );
	NAND3X1 NAND3X1_3549 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_5_), .B(_17376__bF_buf0), .C(_17371__bF_buf3), .Y(_17689_) );
	NAND2X1 NAND2X1_3401 ( .gnd(gnd), .vdd(vdd), .A(_17688_), .B(_17689_), .Y(_17690_) );
	INVX1 INVX1_2238 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_5_), .Y(_17691_) );
	INVX1 INVX1_2239 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_5_), .Y(_17692_) );
	OAI22X1 OAI22X1_192 ( .gnd(gnd), .vdd(vdd), .A(_17691_), .B(_17384__bF_buf4), .C(_17692_), .D(_17383__bF_buf4), .Y(_17693_) );
	NOR2X1 NOR2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_17690_), .B(_17693_), .Y(_17694_) );
	INVX1 INVX1_2240 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_5_), .Y(_17695_) );
	INVX1 INVX1_2241 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_5_), .Y(_17696_) );
	OAI22X1 OAI22X1_193 ( .gnd(gnd), .vdd(vdd), .A(_17695_), .B(_17394__bF_buf4), .C(_17696_), .D(_17393__bF_buf4), .Y(_17697_) );
	INVX1 INVX1_2242 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_5_), .Y(_17698_) );
	INVX1 INVX1_2243 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_5_), .Y(_17699_) );
	OAI22X1 OAI22X1_194 ( .gnd(gnd), .vdd(vdd), .A(_17698_), .B(_17401__bF_buf4), .C(_17699_), .D(_17400__bF_buf4), .Y(_17700_) );
	NOR2X1 NOR2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_17700_), .B(_17697_), .Y(_17701_) );
	NAND2X1 NAND2X1_3402 ( .gnd(gnd), .vdd(vdd), .A(_17694_), .B(_17701_), .Y(_17702_) );
	INVX1 INVX1_2244 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_5_), .Y(_17703_) );
	INVX1 INVX1_2245 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_5_), .Y(_17704_) );
	OAI22X1 OAI22X1_195 ( .gnd(gnd), .vdd(vdd), .A(_17704_), .B(_17408__bF_buf4), .C(_17703_), .D(_17407__bF_buf4), .Y(_17705_) );
	INVX1 INVX1_2246 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_5_), .Y(_17706_) );
	NAND3X1 NAND3X1_3550 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_5_), .B(_17411__bF_buf2), .C(_17413__bF_buf5), .Y(_17707_) );
	OAI21X1 OAI21X1_3562 ( .gnd(gnd), .vdd(vdd), .A(_17706_), .B(_17412__bF_buf4), .C(_17707_), .Y(_17708_) );
	NOR2X1 NOR2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_17705_), .B(_17708_), .Y(_17709_) );
	INVX1 INVX1_2247 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_5_), .Y(_17710_) );
	NAND3X1 NAND3X1_3551 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(registers_r31_5_), .C(_17419__bF_buf4), .Y(_17711_) );
	OAI21X1 OAI21X1_3563 ( .gnd(gnd), .vdd(vdd), .A(_17710_), .B(_17418__bF_buf4), .C(_17711_), .Y(_17712_) );
	INVX1 INVX1_2248 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_5_), .Y(_17713_) );
	NAND3X1 NAND3X1_3552 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_5_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_17714_) );
	OAI21X1 OAI21X1_3564 ( .gnd(gnd), .vdd(vdd), .A(_17713_), .B(_17423__bF_buf4), .C(_17714_), .Y(_17715_) );
	NOR2X1 NOR2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_17712_), .B(_17715_), .Y(_17716_) );
	NAND2X1 NAND2X1_3403 ( .gnd(gnd), .vdd(vdd), .A(_17716_), .B(_17709_), .Y(_17717_) );
	NOR2X1 NOR2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_17717_), .B(_17702_), .Y(_17718_) );
	AOI22X1 AOI22X1_388 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_5_), .C(registers_r1_5_), .D(_17431__bF_buf4), .Y(_17719_) );
	AOI22X1 AOI22X1_389 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_5_), .C(registers_r5_5_), .D(_17436__bF_buf4), .Y(_17720_) );
	INVX1 INVX1_2249 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_5_), .Y(_17721_) );
	NAND3X1 NAND3X1_3553 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_5_), .B(_17432__bF_buf2), .C(_17392__bF_buf7), .Y(_17722_) );
	OAI21X1 OAI21X1_3565 ( .gnd(gnd), .vdd(vdd), .A(_17721_), .B(_17443__bF_buf4), .C(_17722_), .Y(_17723_) );
	AOI21X1 AOI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_5_), .B(_17440__bF_buf4), .C(_17723_), .Y(_17724_) );
	NAND3X1 NAND3X1_3554 ( .gnd(gnd), .vdd(vdd), .A(_17719_), .B(_17720_), .C(_17724_), .Y(_17725_) );
	INVX1 INVX1_2250 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_5_), .Y(_17726_) );
	INVX1 INVX1_2251 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_5_), .Y(_17727_) );
	OAI22X1 OAI22X1_196 ( .gnd(gnd), .vdd(vdd), .A(_17727_), .B(_17450__bF_buf4), .C(_17726_), .D(_17449__bF_buf4), .Y(_17728_) );
	INVX1 INVX1_2252 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_5_), .Y(_17729_) );
	INVX1 INVX1_2253 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_5_), .Y(_17730_) );
	OAI22X1 OAI22X1_197 ( .gnd(gnd), .vdd(vdd), .A(_17729_), .B(_17456__bF_buf4), .C(_17730_), .D(_17454__bF_buf4), .Y(_17731_) );
	NOR2X1 NOR2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_17731_), .B(_17728_), .Y(_17732_) );
	INVX1 INVX1_2254 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_5_), .Y(_17733_) );
	INVX1 INVX1_2255 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_5_), .Y(_17734_) );
	OAI22X1 OAI22X1_198 ( .gnd(gnd), .vdd(vdd), .A(_17733_), .B(_17461__bF_buf4), .C(_17734_), .D(_17462__bF_buf4), .Y(_17735_) );
	INVX1 INVX1_2256 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_5_), .Y(_17736_) );
	INVX1 INVX1_2257 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_5_), .Y(_17737_) );
	OAI22X1 OAI22X1_199 ( .gnd(gnd), .vdd(vdd), .A(_17737_), .B(_17467__bF_buf4), .C(_17736_), .D(_17466__bF_buf4), .Y(_17738_) );
	NOR2X1 NOR2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_17735_), .B(_17738_), .Y(_17739_) );
	NAND2X1 NAND2X1_3404 ( .gnd(gnd), .vdd(vdd), .A(_17732_), .B(_17739_), .Y(_17740_) );
	NOR2X1 NOR2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_17725_), .B(_17740_), .Y(_17741_) );
	NAND2X1 NAND2X1_3405 ( .gnd(gnd), .vdd(vdd), .A(_17741_), .B(_17718_), .Y(_428__5_) );
	NAND3X1 NAND3X1_3555 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_6_), .B(_17373__bF_buf5), .C(_17371__bF_buf2), .Y(_17742_) );
	NAND3X1 NAND3X1_3556 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_6_), .B(_17376__bF_buf5), .C(_17371__bF_buf1), .Y(_17743_) );
	NAND2X1 NAND2X1_3406 ( .gnd(gnd), .vdd(vdd), .A(_17742_), .B(_17743_), .Y(_17744_) );
	INVX1 INVX1_2258 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_6_), .Y(_17745_) );
	INVX1 INVX1_2259 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_6_), .Y(_17746_) );
	OAI22X1 OAI22X1_200 ( .gnd(gnd), .vdd(vdd), .A(_17745_), .B(_17384__bF_buf3), .C(_17746_), .D(_17383__bF_buf3), .Y(_17747_) );
	NOR2X1 NOR2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_17744_), .B(_17747_), .Y(_17748_) );
	INVX1 INVX1_2260 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_6_), .Y(_17749_) );
	INVX1 INVX1_2261 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_6_), .Y(_17750_) );
	OAI22X1 OAI22X1_201 ( .gnd(gnd), .vdd(vdd), .A(_17749_), .B(_17394__bF_buf3), .C(_17750_), .D(_17393__bF_buf3), .Y(_17751_) );
	INVX1 INVX1_2262 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_6_), .Y(_17752_) );
	INVX1 INVX1_2263 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_6_), .Y(_17753_) );
	OAI22X1 OAI22X1_202 ( .gnd(gnd), .vdd(vdd), .A(_17752_), .B(_17401__bF_buf3), .C(_17753_), .D(_17400__bF_buf3), .Y(_17754_) );
	NOR2X1 NOR2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_17754_), .B(_17751_), .Y(_17755_) );
	NAND2X1 NAND2X1_3407 ( .gnd(gnd), .vdd(vdd), .A(_17748_), .B(_17755_), .Y(_17756_) );
	INVX1 INVX1_2264 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_6_), .Y(_17757_) );
	INVX1 INVX1_2265 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_6_), .Y(_17758_) );
	OAI22X1 OAI22X1_203 ( .gnd(gnd), .vdd(vdd), .A(_17758_), .B(_17408__bF_buf3), .C(_17757_), .D(_17407__bF_buf3), .Y(_17759_) );
	INVX1 INVX1_2266 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_6_), .Y(_17760_) );
	NAND3X1 NAND3X1_3557 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_6_), .B(_17411__bF_buf1), .C(_17413__bF_buf3), .Y(_17761_) );
	OAI21X1 OAI21X1_3566 ( .gnd(gnd), .vdd(vdd), .A(_17760_), .B(_17412__bF_buf3), .C(_17761_), .Y(_17762_) );
	NOR2X1 NOR2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_17759_), .B(_17762_), .Y(_17763_) );
	INVX1 INVX1_2267 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_6_), .Y(_17764_) );
	NAND3X1 NAND3X1_3558 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(registers_r31_6_), .C(_17419__bF_buf3), .Y(_17765_) );
	OAI21X1 OAI21X1_3567 ( .gnd(gnd), .vdd(vdd), .A(_17764_), .B(_17418__bF_buf3), .C(_17765_), .Y(_17766_) );
	INVX1 INVX1_2268 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_6_), .Y(_17767_) );
	NAND3X1 NAND3X1_3559 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_6_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_17768_) );
	OAI21X1 OAI21X1_3568 ( .gnd(gnd), .vdd(vdd), .A(_17767_), .B(_17423__bF_buf3), .C(_17768_), .Y(_17769_) );
	NOR2X1 NOR2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_17766_), .B(_17769_), .Y(_17770_) );
	NAND2X1 NAND2X1_3408 ( .gnd(gnd), .vdd(vdd), .A(_17770_), .B(_17763_), .Y(_17771_) );
	NOR2X1 NOR2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_17771_), .B(_17756_), .Y(_17772_) );
	AOI22X1 AOI22X1_390 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_6_), .C(registers_r1_6_), .D(_17431__bF_buf3), .Y(_17773_) );
	AOI22X1 AOI22X1_391 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_6_), .C(registers_r5_6_), .D(_17436__bF_buf3), .Y(_17774_) );
	INVX1 INVX1_2269 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_6_), .Y(_17775_) );
	NAND3X1 NAND3X1_3560 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_6_), .B(_17432__bF_buf1), .C(_17392__bF_buf5), .Y(_17776_) );
	OAI21X1 OAI21X1_3569 ( .gnd(gnd), .vdd(vdd), .A(_17775_), .B(_17443__bF_buf3), .C(_17776_), .Y(_17777_) );
	AOI21X1 AOI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_6_), .B(_17440__bF_buf3), .C(_17777_), .Y(_17778_) );
	NAND3X1 NAND3X1_3561 ( .gnd(gnd), .vdd(vdd), .A(_17773_), .B(_17774_), .C(_17778_), .Y(_17779_) );
	INVX1 INVX1_2270 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_6_), .Y(_17780_) );
	INVX1 INVX1_2271 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_6_), .Y(_17781_) );
	OAI22X1 OAI22X1_204 ( .gnd(gnd), .vdd(vdd), .A(_17781_), .B(_17450__bF_buf3), .C(_17780_), .D(_17449__bF_buf3), .Y(_17782_) );
	INVX1 INVX1_2272 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_6_), .Y(_17783_) );
	INVX1 INVX1_2273 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_6_), .Y(_17784_) );
	OAI22X1 OAI22X1_205 ( .gnd(gnd), .vdd(vdd), .A(_17783_), .B(_17456__bF_buf3), .C(_17784_), .D(_17454__bF_buf3), .Y(_17785_) );
	NOR2X1 NOR2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_17785_), .B(_17782_), .Y(_17786_) );
	INVX1 INVX1_2274 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_6_), .Y(_17787_) );
	INVX1 INVX1_2275 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_6_), .Y(_17788_) );
	OAI22X1 OAI22X1_206 ( .gnd(gnd), .vdd(vdd), .A(_17787_), .B(_17461__bF_buf3), .C(_17788_), .D(_17462__bF_buf3), .Y(_17789_) );
	INVX1 INVX1_2276 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_6_), .Y(_17790_) );
	INVX1 INVX1_2277 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_6_), .Y(_17791_) );
	OAI22X1 OAI22X1_207 ( .gnd(gnd), .vdd(vdd), .A(_17791_), .B(_17467__bF_buf3), .C(_17790_), .D(_17466__bF_buf3), .Y(_17792_) );
	NOR2X1 NOR2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_17789_), .B(_17792_), .Y(_17793_) );
	NAND2X1 NAND2X1_3409 ( .gnd(gnd), .vdd(vdd), .A(_17786_), .B(_17793_), .Y(_17794_) );
	NOR2X1 NOR2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_17779_), .B(_17794_), .Y(_17795_) );
	NAND2X1 NAND2X1_3410 ( .gnd(gnd), .vdd(vdd), .A(_17795_), .B(_17772_), .Y(_428__6_) );
	NAND3X1 NAND3X1_3562 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_7_), .B(_17373__bF_buf4), .C(_17371__bF_buf0), .Y(_17796_) );
	NAND3X1 NAND3X1_3563 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_7_), .B(_17376__bF_buf4), .C(_17371__bF_buf7), .Y(_17797_) );
	NAND2X1 NAND2X1_3411 ( .gnd(gnd), .vdd(vdd), .A(_17796_), .B(_17797_), .Y(_17798_) );
	INVX1 INVX1_2278 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_7_), .Y(_17799_) );
	INVX1 INVX1_2279 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_7_), .Y(_17800_) );
	OAI22X1 OAI22X1_208 ( .gnd(gnd), .vdd(vdd), .A(_17799_), .B(_17384__bF_buf2), .C(_17800_), .D(_17383__bF_buf2), .Y(_17801_) );
	NOR2X1 NOR2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_17798_), .B(_17801_), .Y(_17802_) );
	INVX1 INVX1_2280 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_7_), .Y(_17803_) );
	INVX1 INVX1_2281 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_7_), .Y(_17804_) );
	OAI22X1 OAI22X1_209 ( .gnd(gnd), .vdd(vdd), .A(_17803_), .B(_17394__bF_buf2), .C(_17804_), .D(_17393__bF_buf2), .Y(_17805_) );
	INVX1 INVX1_2282 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_7_), .Y(_17806_) );
	INVX1 INVX1_2283 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_7_), .Y(_17807_) );
	OAI22X1 OAI22X1_210 ( .gnd(gnd), .vdd(vdd), .A(_17806_), .B(_17401__bF_buf2), .C(_17807_), .D(_17400__bF_buf2), .Y(_17808_) );
	NOR2X1 NOR2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_17808_), .B(_17805_), .Y(_17809_) );
	NAND2X1 NAND2X1_3412 ( .gnd(gnd), .vdd(vdd), .A(_17802_), .B(_17809_), .Y(_17810_) );
	INVX1 INVX1_2284 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_7_), .Y(_17811_) );
	INVX1 INVX1_2285 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_7_), .Y(_17812_) );
	OAI22X1 OAI22X1_211 ( .gnd(gnd), .vdd(vdd), .A(_17812_), .B(_17408__bF_buf2), .C(_17811_), .D(_17407__bF_buf2), .Y(_17813_) );
	INVX1 INVX1_2286 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_7_), .Y(_17814_) );
	NAND3X1 NAND3X1_3564 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_7_), .B(_17411__bF_buf0), .C(_17413__bF_buf1), .Y(_17815_) );
	OAI21X1 OAI21X1_3570 ( .gnd(gnd), .vdd(vdd), .A(_17814_), .B(_17412__bF_buf2), .C(_17815_), .Y(_17816_) );
	NOR2X1 NOR2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_17813_), .B(_17816_), .Y(_17817_) );
	INVX1 INVX1_2287 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_7_), .Y(_17818_) );
	NAND3X1 NAND3X1_3565 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(registers_r31_7_), .C(_17419__bF_buf2), .Y(_17819_) );
	OAI21X1 OAI21X1_3571 ( .gnd(gnd), .vdd(vdd), .A(_17818_), .B(_17418__bF_buf2), .C(_17819_), .Y(_17820_) );
	INVX1 INVX1_2288 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_7_), .Y(_17821_) );
	NAND3X1 NAND3X1_3566 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_7_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_17822_) );
	OAI21X1 OAI21X1_3572 ( .gnd(gnd), .vdd(vdd), .A(_17821_), .B(_17423__bF_buf2), .C(_17822_), .Y(_17823_) );
	NOR2X1 NOR2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_17820_), .B(_17823_), .Y(_17824_) );
	NAND2X1 NAND2X1_3413 ( .gnd(gnd), .vdd(vdd), .A(_17824_), .B(_17817_), .Y(_17825_) );
	NOR2X1 NOR2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_17825_), .B(_17810_), .Y(_17826_) );
	AOI22X1 AOI22X1_392 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf2), .B(registers_a2_7_), .C(registers_r1_7_), .D(_17431__bF_buf2), .Y(_17827_) );
	AOI22X1 AOI22X1_393 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf2), .B(registers_r4_7_), .C(registers_r5_7_), .D(_17436__bF_buf2), .Y(_17828_) );
	INVX1 INVX1_2289 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_7_), .Y(_17829_) );
	NAND3X1 NAND3X1_3567 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_7_), .B(_17432__bF_buf0), .C(_17392__bF_buf3), .Y(_17830_) );
	OAI21X1 OAI21X1_3573 ( .gnd(gnd), .vdd(vdd), .A(_17829_), .B(_17443__bF_buf2), .C(_17830_), .Y(_17831_) );
	AOI21X1 AOI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_7_), .B(_17440__bF_buf2), .C(_17831_), .Y(_17832_) );
	NAND3X1 NAND3X1_3568 ( .gnd(gnd), .vdd(vdd), .A(_17827_), .B(_17828_), .C(_17832_), .Y(_17833_) );
	INVX1 INVX1_2290 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_7_), .Y(_17834_) );
	INVX1 INVX1_2291 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_7_), .Y(_17835_) );
	OAI22X1 OAI22X1_212 ( .gnd(gnd), .vdd(vdd), .A(_17835_), .B(_17450__bF_buf2), .C(_17834_), .D(_17449__bF_buf2), .Y(_17836_) );
	INVX1 INVX1_2292 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_7_), .Y(_17837_) );
	INVX1 INVX1_2293 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_7_), .Y(_17838_) );
	OAI22X1 OAI22X1_213 ( .gnd(gnd), .vdd(vdd), .A(_17837_), .B(_17456__bF_buf2), .C(_17838_), .D(_17454__bF_buf2), .Y(_17839_) );
	NOR2X1 NOR2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_17839_), .B(_17836_), .Y(_17840_) );
	INVX1 INVX1_2294 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_7_), .Y(_17841_) );
	INVX1 INVX1_2295 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_7_), .Y(_17842_) );
	OAI22X1 OAI22X1_214 ( .gnd(gnd), .vdd(vdd), .A(_17841_), .B(_17461__bF_buf2), .C(_17842_), .D(_17462__bF_buf2), .Y(_17843_) );
	INVX1 INVX1_2296 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_7_), .Y(_17844_) );
	INVX1 INVX1_2297 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_7_), .Y(_17845_) );
	OAI22X1 OAI22X1_215 ( .gnd(gnd), .vdd(vdd), .A(_17845_), .B(_17467__bF_buf2), .C(_17844_), .D(_17466__bF_buf2), .Y(_17846_) );
	NOR2X1 NOR2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_17843_), .B(_17846_), .Y(_17847_) );
	NAND2X1 NAND2X1_3414 ( .gnd(gnd), .vdd(vdd), .A(_17840_), .B(_17847_), .Y(_17848_) );
	NOR2X1 NOR2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_17833_), .B(_17848_), .Y(_17849_) );
	NAND2X1 NAND2X1_3415 ( .gnd(gnd), .vdd(vdd), .A(_17849_), .B(_17826_), .Y(_428__7_) );
	NAND3X1 NAND3X1_3569 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_8_), .B(_17373__bF_buf3), .C(_17371__bF_buf6), .Y(_17850_) );
	NAND3X1 NAND3X1_3570 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_8_), .B(_17376__bF_buf3), .C(_17371__bF_buf5), .Y(_17851_) );
	NAND2X1 NAND2X1_3416 ( .gnd(gnd), .vdd(vdd), .A(_17850_), .B(_17851_), .Y(_17852_) );
	INVX1 INVX1_2298 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_8_), .Y(_17853_) );
	INVX1 INVX1_2299 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_8_), .Y(_17854_) );
	OAI22X1 OAI22X1_216 ( .gnd(gnd), .vdd(vdd), .A(_17853_), .B(_17384__bF_buf1), .C(_17854_), .D(_17383__bF_buf1), .Y(_17855_) );
	NOR2X1 NOR2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_17852_), .B(_17855_), .Y(_17856_) );
	INVX1 INVX1_2300 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_8_), .Y(_17857_) );
	INVX1 INVX1_2301 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_8_), .Y(_17858_) );
	OAI22X1 OAI22X1_217 ( .gnd(gnd), .vdd(vdd), .A(_17857_), .B(_17394__bF_buf1), .C(_17858_), .D(_17393__bF_buf1), .Y(_17859_) );
	INVX1 INVX1_2302 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_8_), .Y(_17860_) );
	INVX1 INVX1_2303 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_8_), .Y(_17861_) );
	OAI22X1 OAI22X1_218 ( .gnd(gnd), .vdd(vdd), .A(_17860_), .B(_17401__bF_buf1), .C(_17861_), .D(_17400__bF_buf1), .Y(_17862_) );
	NOR2X1 NOR2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_17862_), .B(_17859_), .Y(_17863_) );
	NAND2X1 NAND2X1_3417 ( .gnd(gnd), .vdd(vdd), .A(_17856_), .B(_17863_), .Y(_17864_) );
	INVX1 INVX1_2304 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_8_), .Y(_17865_) );
	INVX1 INVX1_2305 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_8_), .Y(_17866_) );
	OAI22X1 OAI22X1_219 ( .gnd(gnd), .vdd(vdd), .A(_17866_), .B(_17408__bF_buf1), .C(_17865_), .D(_17407__bF_buf1), .Y(_17867_) );
	INVX1 INVX1_2306 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_8_), .Y(_17868_) );
	NAND3X1 NAND3X1_3571 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_8_), .B(_17411__bF_buf5), .C(_17413__bF_buf7), .Y(_17869_) );
	OAI21X1 OAI21X1_3574 ( .gnd(gnd), .vdd(vdd), .A(_17868_), .B(_17412__bF_buf1), .C(_17869_), .Y(_17870_) );
	NOR2X1 NOR2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_17867_), .B(_17870_), .Y(_17871_) );
	INVX1 INVX1_2307 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_8_), .Y(_17872_) );
	NAND3X1 NAND3X1_3572 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(registers_r31_8_), .C(_17419__bF_buf1), .Y(_17873_) );
	OAI21X1 OAI21X1_3575 ( .gnd(gnd), .vdd(vdd), .A(_17872_), .B(_17418__bF_buf1), .C(_17873_), .Y(_17874_) );
	INVX1 INVX1_2308 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_8_), .Y(_17875_) );
	NAND3X1 NAND3X1_3573 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_8_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_17876_) );
	OAI21X1 OAI21X1_3576 ( .gnd(gnd), .vdd(vdd), .A(_17875_), .B(_17423__bF_buf1), .C(_17876_), .Y(_17877_) );
	NOR2X1 NOR2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_17874_), .B(_17877_), .Y(_17878_) );
	NAND2X1 NAND2X1_3418 ( .gnd(gnd), .vdd(vdd), .A(_17878_), .B(_17871_), .Y(_17879_) );
	NOR2X1 NOR2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_17879_), .B(_17864_), .Y(_17880_) );
	AOI22X1 AOI22X1_394 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf1), .B(registers_a2_8_), .C(registers_r1_8_), .D(_17431__bF_buf1), .Y(_17881_) );
	AOI22X1 AOI22X1_395 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf1), .B(registers_r4_8_), .C(registers_r5_8_), .D(_17436__bF_buf1), .Y(_17882_) );
	INVX1 INVX1_2309 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_8_), .Y(_17883_) );
	NAND3X1 NAND3X1_3574 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_8_), .B(_17432__bF_buf4), .C(_17392__bF_buf1), .Y(_17884_) );
	OAI21X1 OAI21X1_3577 ( .gnd(gnd), .vdd(vdd), .A(_17883_), .B(_17443__bF_buf1), .C(_17884_), .Y(_17885_) );
	AOI21X1 AOI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_8_), .B(_17440__bF_buf1), .C(_17885_), .Y(_17886_) );
	NAND3X1 NAND3X1_3575 ( .gnd(gnd), .vdd(vdd), .A(_17881_), .B(_17882_), .C(_17886_), .Y(_17887_) );
	INVX1 INVX1_2310 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_8_), .Y(_17888_) );
	INVX1 INVX1_2311 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_8_), .Y(_17889_) );
	OAI22X1 OAI22X1_220 ( .gnd(gnd), .vdd(vdd), .A(_17889_), .B(_17450__bF_buf1), .C(_17888_), .D(_17449__bF_buf1), .Y(_17890_) );
	INVX1 INVX1_2312 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_8_), .Y(_17891_) );
	INVX1 INVX1_2313 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_8_), .Y(_17892_) );
	OAI22X1 OAI22X1_221 ( .gnd(gnd), .vdd(vdd), .A(_17891_), .B(_17456__bF_buf1), .C(_17892_), .D(_17454__bF_buf1), .Y(_17893_) );
	NOR2X1 NOR2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_17893_), .B(_17890_), .Y(_17894_) );
	INVX1 INVX1_2314 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_8_), .Y(_17895_) );
	INVX1 INVX1_2315 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_8_), .Y(_17896_) );
	OAI22X1 OAI22X1_222 ( .gnd(gnd), .vdd(vdd), .A(_17895_), .B(_17461__bF_buf1), .C(_17896_), .D(_17462__bF_buf1), .Y(_17897_) );
	INVX1 INVX1_2316 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_8_), .Y(_17898_) );
	INVX1 INVX1_2317 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_8_), .Y(_17899_) );
	OAI22X1 OAI22X1_223 ( .gnd(gnd), .vdd(vdd), .A(_17899_), .B(_17467__bF_buf1), .C(_17898_), .D(_17466__bF_buf1), .Y(_17900_) );
	NOR2X1 NOR2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_17897_), .B(_17900_), .Y(_17901_) );
	NAND2X1 NAND2X1_3419 ( .gnd(gnd), .vdd(vdd), .A(_17894_), .B(_17901_), .Y(_17902_) );
	NOR2X1 NOR2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_17887_), .B(_17902_), .Y(_17903_) );
	NAND2X1 NAND2X1_3420 ( .gnd(gnd), .vdd(vdd), .A(_17903_), .B(_17880_), .Y(_428__8_) );
	NAND3X1 NAND3X1_3576 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_9_), .B(_17373__bF_buf2), .C(_17371__bF_buf4), .Y(_17904_) );
	NAND3X1 NAND3X1_3577 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_9_), .B(_17376__bF_buf2), .C(_17371__bF_buf3), .Y(_17905_) );
	NAND2X1 NAND2X1_3421 ( .gnd(gnd), .vdd(vdd), .A(_17904_), .B(_17905_), .Y(_17906_) );
	INVX1 INVX1_2318 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_9_), .Y(_17907_) );
	INVX1 INVX1_2319 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_9_), .Y(_17908_) );
	OAI22X1 OAI22X1_224 ( .gnd(gnd), .vdd(vdd), .A(_17907_), .B(_17384__bF_buf0), .C(_17908_), .D(_17383__bF_buf0), .Y(_17909_) );
	NOR2X1 NOR2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_17906_), .B(_17909_), .Y(_17910_) );
	INVX1 INVX1_2320 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_9_), .Y(_17911_) );
	INVX1 INVX1_2321 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_9_), .Y(_17912_) );
	OAI22X1 OAI22X1_225 ( .gnd(gnd), .vdd(vdd), .A(_17911_), .B(_17394__bF_buf0), .C(_17912_), .D(_17393__bF_buf0), .Y(_17913_) );
	INVX1 INVX1_2322 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_9_), .Y(_17914_) );
	INVX1 INVX1_2323 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_9_), .Y(_17915_) );
	OAI22X1 OAI22X1_226 ( .gnd(gnd), .vdd(vdd), .A(_17914_), .B(_17401__bF_buf0), .C(_17915_), .D(_17400__bF_buf0), .Y(_17916_) );
	NOR2X1 NOR2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_17916_), .B(_17913_), .Y(_17917_) );
	NAND2X1 NAND2X1_3422 ( .gnd(gnd), .vdd(vdd), .A(_17910_), .B(_17917_), .Y(_17918_) );
	INVX1 INVX1_2324 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_9_), .Y(_17919_) );
	INVX1 INVX1_2325 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_9_), .Y(_17920_) );
	OAI22X1 OAI22X1_227 ( .gnd(gnd), .vdd(vdd), .A(_17920_), .B(_17408__bF_buf0), .C(_17919_), .D(_17407__bF_buf0), .Y(_17921_) );
	INVX1 INVX1_2326 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_9_), .Y(_17922_) );
	NAND3X1 NAND3X1_3578 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_9_), .B(_17411__bF_buf4), .C(_17413__bF_buf5), .Y(_17923_) );
	OAI21X1 OAI21X1_3578 ( .gnd(gnd), .vdd(vdd), .A(_17922_), .B(_17412__bF_buf0), .C(_17923_), .Y(_17924_) );
	NOR2X1 NOR2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_17921_), .B(_17924_), .Y(_17925_) );
	INVX1 INVX1_2327 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_9_), .Y(_17926_) );
	NAND3X1 NAND3X1_3579 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(registers_r31_9_), .C(_17419__bF_buf0), .Y(_17927_) );
	OAI21X1 OAI21X1_3579 ( .gnd(gnd), .vdd(vdd), .A(_17926_), .B(_17418__bF_buf0), .C(_17927_), .Y(_17928_) );
	INVX1 INVX1_2328 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_9_), .Y(_17929_) );
	NAND3X1 NAND3X1_3580 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_9_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_17930_) );
	OAI21X1 OAI21X1_3580 ( .gnd(gnd), .vdd(vdd), .A(_17929_), .B(_17423__bF_buf0), .C(_17930_), .Y(_17931_) );
	NOR2X1 NOR2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_17928_), .B(_17931_), .Y(_17932_) );
	NAND2X1 NAND2X1_3423 ( .gnd(gnd), .vdd(vdd), .A(_17932_), .B(_17925_), .Y(_17933_) );
	NOR2X1 NOR2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_17933_), .B(_17918_), .Y(_17934_) );
	AOI22X1 AOI22X1_396 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf0), .B(registers_a2_9_), .C(registers_r1_9_), .D(_17431__bF_buf0), .Y(_17935_) );
	AOI22X1 AOI22X1_397 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf0), .B(registers_r4_9_), .C(registers_r5_9_), .D(_17436__bF_buf0), .Y(_17936_) );
	INVX1 INVX1_2329 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_9_), .Y(_17937_) );
	NAND3X1 NAND3X1_3581 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_9_), .B(_17432__bF_buf3), .C(_17392__bF_buf7), .Y(_17938_) );
	OAI21X1 OAI21X1_3581 ( .gnd(gnd), .vdd(vdd), .A(_17937_), .B(_17443__bF_buf0), .C(_17938_), .Y(_17939_) );
	AOI21X1 AOI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_9_), .B(_17440__bF_buf0), .C(_17939_), .Y(_17940_) );
	NAND3X1 NAND3X1_3582 ( .gnd(gnd), .vdd(vdd), .A(_17935_), .B(_17936_), .C(_17940_), .Y(_17941_) );
	INVX1 INVX1_2330 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_9_), .Y(_17942_) );
	INVX1 INVX1_2331 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_9_), .Y(_17943_) );
	OAI22X1 OAI22X1_228 ( .gnd(gnd), .vdd(vdd), .A(_17943_), .B(_17450__bF_buf0), .C(_17942_), .D(_17449__bF_buf0), .Y(_17944_) );
	INVX1 INVX1_2332 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_9_), .Y(_17945_) );
	INVX1 INVX1_2333 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_9_), .Y(_17946_) );
	OAI22X1 OAI22X1_229 ( .gnd(gnd), .vdd(vdd), .A(_17945_), .B(_17456__bF_buf0), .C(_17946_), .D(_17454__bF_buf0), .Y(_17947_) );
	NOR2X1 NOR2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_17947_), .B(_17944_), .Y(_17948_) );
	INVX1 INVX1_2334 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_9_), .Y(_17949_) );
	INVX1 INVX1_2335 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_9_), .Y(_17950_) );
	OAI22X1 OAI22X1_230 ( .gnd(gnd), .vdd(vdd), .A(_17949_), .B(_17461__bF_buf0), .C(_17950_), .D(_17462__bF_buf0), .Y(_17951_) );
	INVX1 INVX1_2336 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_9_), .Y(_17952_) );
	INVX1 INVX1_2337 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_9_), .Y(_17953_) );
	OAI22X1 OAI22X1_231 ( .gnd(gnd), .vdd(vdd), .A(_17953_), .B(_17467__bF_buf0), .C(_17952_), .D(_17466__bF_buf0), .Y(_17954_) );
	NOR2X1 NOR2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_17951_), .B(_17954_), .Y(_17955_) );
	NAND2X1 NAND2X1_3424 ( .gnd(gnd), .vdd(vdd), .A(_17948_), .B(_17955_), .Y(_17956_) );
	NOR2X1 NOR2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_17941_), .B(_17956_), .Y(_17957_) );
	NAND2X1 NAND2X1_3425 ( .gnd(gnd), .vdd(vdd), .A(_17957_), .B(_17934_), .Y(_428__9_) );
	NAND3X1 NAND3X1_3583 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_10_), .B(_17373__bF_buf1), .C(_17371__bF_buf2), .Y(_17958_) );
	NAND3X1 NAND3X1_3584 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_10_), .B(_17376__bF_buf1), .C(_17371__bF_buf1), .Y(_17959_) );
	NAND2X1 NAND2X1_3426 ( .gnd(gnd), .vdd(vdd), .A(_17958_), .B(_17959_), .Y(_17960_) );
	INVX1 INVX1_2338 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_10_), .Y(_17961_) );
	INVX1 INVX1_2339 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_10_), .Y(_17962_) );
	OAI22X1 OAI22X1_232 ( .gnd(gnd), .vdd(vdd), .A(_17961_), .B(_17384__bF_buf4), .C(_17962_), .D(_17383__bF_buf4), .Y(_17963_) );
	NOR2X1 NOR2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_17960_), .B(_17963_), .Y(_17964_) );
	INVX1 INVX1_2340 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_10_), .Y(_17965_) );
	INVX1 INVX1_2341 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_10_), .Y(_17966_) );
	OAI22X1 OAI22X1_233 ( .gnd(gnd), .vdd(vdd), .A(_17965_), .B(_17394__bF_buf4), .C(_17966_), .D(_17393__bF_buf4), .Y(_17967_) );
	INVX1 INVX1_2342 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_10_), .Y(_17968_) );
	INVX1 INVX1_2343 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_10_), .Y(_17969_) );
	OAI22X1 OAI22X1_234 ( .gnd(gnd), .vdd(vdd), .A(_17968_), .B(_17401__bF_buf4), .C(_17969_), .D(_17400__bF_buf4), .Y(_17970_) );
	NOR2X1 NOR2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_17970_), .B(_17967_), .Y(_17971_) );
	NAND2X1 NAND2X1_3427 ( .gnd(gnd), .vdd(vdd), .A(_17964_), .B(_17971_), .Y(_17972_) );
	INVX1 INVX1_2344 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_10_), .Y(_17973_) );
	INVX1 INVX1_2345 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_10_), .Y(_17974_) );
	OAI22X1 OAI22X1_235 ( .gnd(gnd), .vdd(vdd), .A(_17974_), .B(_17408__bF_buf4), .C(_17973_), .D(_17407__bF_buf4), .Y(_17975_) );
	INVX1 INVX1_2346 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_10_), .Y(_17976_) );
	NAND3X1 NAND3X1_3585 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_10_), .B(_17411__bF_buf3), .C(_17413__bF_buf3), .Y(_17977_) );
	OAI21X1 OAI21X1_3582 ( .gnd(gnd), .vdd(vdd), .A(_17976_), .B(_17412__bF_buf4), .C(_17977_), .Y(_17978_) );
	NOR2X1 NOR2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_17975_), .B(_17978_), .Y(_17979_) );
	INVX1 INVX1_2347 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_10_), .Y(_17980_) );
	NAND3X1 NAND3X1_3586 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(registers_r31_10_), .C(_17419__bF_buf4), .Y(_17981_) );
	OAI21X1 OAI21X1_3583 ( .gnd(gnd), .vdd(vdd), .A(_17980_), .B(_17418__bF_buf4), .C(_17981_), .Y(_17982_) );
	INVX1 INVX1_2348 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_10_), .Y(_17983_) );
	NAND3X1 NAND3X1_3587 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_10_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_17984_) );
	OAI21X1 OAI21X1_3584 ( .gnd(gnd), .vdd(vdd), .A(_17983_), .B(_17423__bF_buf4), .C(_17984_), .Y(_17985_) );
	NOR2X1 NOR2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_17982_), .B(_17985_), .Y(_17986_) );
	NAND2X1 NAND2X1_3428 ( .gnd(gnd), .vdd(vdd), .A(_17986_), .B(_17979_), .Y(_17987_) );
	NOR2X1 NOR2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_17987_), .B(_17972_), .Y(_17988_) );
	AOI22X1 AOI22X1_398 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_10_), .C(registers_r1_10_), .D(_17431__bF_buf4), .Y(_17989_) );
	AOI22X1 AOI22X1_399 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_10_), .C(registers_r5_10_), .D(_17436__bF_buf4), .Y(_17990_) );
	INVX1 INVX1_2349 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_10_), .Y(_17991_) );
	NAND3X1 NAND3X1_3588 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_10_), .B(_17432__bF_buf2), .C(_17392__bF_buf5), .Y(_17992_) );
	OAI21X1 OAI21X1_3585 ( .gnd(gnd), .vdd(vdd), .A(_17991_), .B(_17443__bF_buf4), .C(_17992_), .Y(_17993_) );
	AOI21X1 AOI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_10_), .B(_17440__bF_buf4), .C(_17993_), .Y(_17994_) );
	NAND3X1 NAND3X1_3589 ( .gnd(gnd), .vdd(vdd), .A(_17989_), .B(_17990_), .C(_17994_), .Y(_17995_) );
	INVX1 INVX1_2350 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_10_), .Y(_17996_) );
	INVX1 INVX1_2351 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_10_), .Y(_17997_) );
	OAI22X1 OAI22X1_236 ( .gnd(gnd), .vdd(vdd), .A(_17997_), .B(_17450__bF_buf4), .C(_17996_), .D(_17449__bF_buf4), .Y(_17998_) );
	INVX1 INVX1_2352 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_10_), .Y(_17999_) );
	INVX1 INVX1_2353 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_10_), .Y(_18000_) );
	OAI22X1 OAI22X1_237 ( .gnd(gnd), .vdd(vdd), .A(_17999_), .B(_17456__bF_buf4), .C(_18000_), .D(_17454__bF_buf4), .Y(_18001_) );
	NOR2X1 NOR2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_18001_), .B(_17998_), .Y(_18002_) );
	INVX1 INVX1_2354 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_10_), .Y(_18003_) );
	INVX1 INVX1_2355 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_10_), .Y(_18004_) );
	OAI22X1 OAI22X1_238 ( .gnd(gnd), .vdd(vdd), .A(_18003_), .B(_17461__bF_buf4), .C(_18004_), .D(_17462__bF_buf4), .Y(_18005_) );
	INVX1 INVX1_2356 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_10_), .Y(_18006_) );
	INVX1 INVX1_2357 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_10_), .Y(_18007_) );
	OAI22X1 OAI22X1_239 ( .gnd(gnd), .vdd(vdd), .A(_18007_), .B(_17467__bF_buf4), .C(_18006_), .D(_17466__bF_buf4), .Y(_18008_) );
	NOR2X1 NOR2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_18005_), .B(_18008_), .Y(_18009_) );
	NAND2X1 NAND2X1_3429 ( .gnd(gnd), .vdd(vdd), .A(_18002_), .B(_18009_), .Y(_18010_) );
	NOR2X1 NOR2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_17995_), .B(_18010_), .Y(_18011_) );
	NAND2X1 NAND2X1_3430 ( .gnd(gnd), .vdd(vdd), .A(_18011_), .B(_17988_), .Y(_428__10_) );
	NAND3X1 NAND3X1_3590 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_11_), .B(_17373__bF_buf0), .C(_17371__bF_buf0), .Y(_18012_) );
	NAND3X1 NAND3X1_3591 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_11_), .B(_17376__bF_buf0), .C(_17371__bF_buf7), .Y(_18013_) );
	NAND2X1 NAND2X1_3431 ( .gnd(gnd), .vdd(vdd), .A(_18012_), .B(_18013_), .Y(_18014_) );
	INVX1 INVX1_2358 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_11_), .Y(_18015_) );
	INVX1 INVX1_2359 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_11_), .Y(_18016_) );
	OAI22X1 OAI22X1_240 ( .gnd(gnd), .vdd(vdd), .A(_18015_), .B(_17384__bF_buf3), .C(_18016_), .D(_17383__bF_buf3), .Y(_18017_) );
	NOR2X1 NOR2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_18014_), .B(_18017_), .Y(_18018_) );
	INVX1 INVX1_2360 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_11_), .Y(_18019_) );
	INVX1 INVX1_2361 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_11_), .Y(_18020_) );
	OAI22X1 OAI22X1_241 ( .gnd(gnd), .vdd(vdd), .A(_18019_), .B(_17394__bF_buf3), .C(_18020_), .D(_17393__bF_buf3), .Y(_18021_) );
	INVX1 INVX1_2362 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_11_), .Y(_18022_) );
	INVX1 INVX1_2363 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_11_), .Y(_18023_) );
	OAI22X1 OAI22X1_242 ( .gnd(gnd), .vdd(vdd), .A(_18022_), .B(_17401__bF_buf3), .C(_18023_), .D(_17400__bF_buf3), .Y(_18024_) );
	NOR2X1 NOR2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_18024_), .B(_18021_), .Y(_18025_) );
	NAND2X1 NAND2X1_3432 ( .gnd(gnd), .vdd(vdd), .A(_18018_), .B(_18025_), .Y(_18026_) );
	INVX1 INVX1_2364 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_11_), .Y(_18027_) );
	INVX1 INVX1_2365 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_11_), .Y(_18028_) );
	OAI22X1 OAI22X1_243 ( .gnd(gnd), .vdd(vdd), .A(_18028_), .B(_17408__bF_buf3), .C(_18027_), .D(_17407__bF_buf3), .Y(_18029_) );
	INVX1 INVX1_2366 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_11_), .Y(_18030_) );
	NAND3X1 NAND3X1_3592 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_11_), .B(_17411__bF_buf2), .C(_17413__bF_buf1), .Y(_18031_) );
	OAI21X1 OAI21X1_3586 ( .gnd(gnd), .vdd(vdd), .A(_18030_), .B(_17412__bF_buf3), .C(_18031_), .Y(_18032_) );
	NOR2X1 NOR2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_18029_), .B(_18032_), .Y(_18033_) );
	INVX1 INVX1_2367 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_11_), .Y(_18034_) );
	NAND3X1 NAND3X1_3593 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .B(registers_r31_11_), .C(_17419__bF_buf3), .Y(_18035_) );
	OAI21X1 OAI21X1_3587 ( .gnd(gnd), .vdd(vdd), .A(_18034_), .B(_17418__bF_buf3), .C(_18035_), .Y(_18036_) );
	INVX1 INVX1_2368 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_11_), .Y(_18037_) );
	NAND3X1 NAND3X1_3594 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_11_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_18038_) );
	OAI21X1 OAI21X1_3588 ( .gnd(gnd), .vdd(vdd), .A(_18037_), .B(_17423__bF_buf3), .C(_18038_), .Y(_18039_) );
	NOR2X1 NOR2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_18036_), .B(_18039_), .Y(_18040_) );
	NAND2X1 NAND2X1_3433 ( .gnd(gnd), .vdd(vdd), .A(_18040_), .B(_18033_), .Y(_18041_) );
	NOR2X1 NOR2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_18041_), .B(_18026_), .Y(_18042_) );
	AOI22X1 AOI22X1_400 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_11_), .C(registers_r1_11_), .D(_17431__bF_buf3), .Y(_18043_) );
	AOI22X1 AOI22X1_401 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_11_), .C(registers_r5_11_), .D(_17436__bF_buf3), .Y(_18044_) );
	INVX1 INVX1_2369 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_11_), .Y(_18045_) );
	NAND3X1 NAND3X1_3595 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_11_), .B(_17432__bF_buf1), .C(_17392__bF_buf3), .Y(_18046_) );
	OAI21X1 OAI21X1_3589 ( .gnd(gnd), .vdd(vdd), .A(_18045_), .B(_17443__bF_buf3), .C(_18046_), .Y(_18047_) );
	AOI21X1 AOI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_11_), .B(_17440__bF_buf3), .C(_18047_), .Y(_18048_) );
	NAND3X1 NAND3X1_3596 ( .gnd(gnd), .vdd(vdd), .A(_18043_), .B(_18044_), .C(_18048_), .Y(_18049_) );
	INVX1 INVX1_2370 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_11_), .Y(_18050_) );
	INVX1 INVX1_2371 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_11_), .Y(_18051_) );
	OAI22X1 OAI22X1_244 ( .gnd(gnd), .vdd(vdd), .A(_18051_), .B(_17450__bF_buf3), .C(_18050_), .D(_17449__bF_buf3), .Y(_18052_) );
	INVX1 INVX1_2372 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_11_), .Y(_18053_) );
	INVX1 INVX1_2373 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_11_), .Y(_18054_) );
	OAI22X1 OAI22X1_245 ( .gnd(gnd), .vdd(vdd), .A(_18053_), .B(_17456__bF_buf3), .C(_18054_), .D(_17454__bF_buf3), .Y(_18055_) );
	NOR2X1 NOR2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_18055_), .B(_18052_), .Y(_18056_) );
	INVX1 INVX1_2374 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_11_), .Y(_18057_) );
	INVX1 INVX1_2375 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_11_), .Y(_18058_) );
	OAI22X1 OAI22X1_246 ( .gnd(gnd), .vdd(vdd), .A(_18057_), .B(_17461__bF_buf3), .C(_18058_), .D(_17462__bF_buf3), .Y(_18059_) );
	INVX1 INVX1_2376 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_11_), .Y(_18060_) );
	INVX1 INVX1_2377 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_11_), .Y(_18061_) );
	OAI22X1 OAI22X1_247 ( .gnd(gnd), .vdd(vdd), .A(_18061_), .B(_17467__bF_buf3), .C(_18060_), .D(_17466__bF_buf3), .Y(_18062_) );
	NOR2X1 NOR2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_18059_), .B(_18062_), .Y(_18063_) );
	NAND2X1 NAND2X1_3434 ( .gnd(gnd), .vdd(vdd), .A(_18056_), .B(_18063_), .Y(_18064_) );
	NOR2X1 NOR2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_18049_), .B(_18064_), .Y(_18065_) );
	NAND2X1 NAND2X1_3435 ( .gnd(gnd), .vdd(vdd), .A(_18065_), .B(_18042_), .Y(_428__11_) );
	NAND3X1 NAND3X1_3597 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_12_), .B(_17373__bF_buf5), .C(_17371__bF_buf6), .Y(_18066_) );
	NAND3X1 NAND3X1_3598 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_12_), .B(_17376__bF_buf5), .C(_17371__bF_buf5), .Y(_18067_) );
	NAND2X1 NAND2X1_3436 ( .gnd(gnd), .vdd(vdd), .A(_18066_), .B(_18067_), .Y(_18068_) );
	INVX1 INVX1_2378 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_12_), .Y(_18069_) );
	INVX1 INVX1_2379 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_12_), .Y(_18070_) );
	OAI22X1 OAI22X1_248 ( .gnd(gnd), .vdd(vdd), .A(_18069_), .B(_17384__bF_buf2), .C(_18070_), .D(_17383__bF_buf2), .Y(_18071_) );
	NOR2X1 NOR2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_18068_), .B(_18071_), .Y(_18072_) );
	INVX1 INVX1_2380 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_12_), .Y(_18073_) );
	INVX1 INVX1_2381 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_12_), .Y(_18074_) );
	OAI22X1 OAI22X1_249 ( .gnd(gnd), .vdd(vdd), .A(_18073_), .B(_17394__bF_buf2), .C(_18074_), .D(_17393__bF_buf2), .Y(_18075_) );
	INVX1 INVX1_2382 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_12_), .Y(_18076_) );
	INVX1 INVX1_2383 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_12_), .Y(_18077_) );
	OAI22X1 OAI22X1_250 ( .gnd(gnd), .vdd(vdd), .A(_18076_), .B(_17401__bF_buf2), .C(_18077_), .D(_17400__bF_buf2), .Y(_18078_) );
	NOR2X1 NOR2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_18078_), .B(_18075_), .Y(_18079_) );
	NAND2X1 NAND2X1_3437 ( .gnd(gnd), .vdd(vdd), .A(_18072_), .B(_18079_), .Y(_18080_) );
	INVX1 INVX1_2384 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_12_), .Y(_18081_) );
	INVX1 INVX1_2385 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_12_), .Y(_18082_) );
	OAI22X1 OAI22X1_251 ( .gnd(gnd), .vdd(vdd), .A(_18082_), .B(_17408__bF_buf2), .C(_18081_), .D(_17407__bF_buf2), .Y(_18083_) );
	INVX1 INVX1_2386 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_12_), .Y(_18084_) );
	NAND3X1 NAND3X1_3599 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_12_), .B(_17411__bF_buf1), .C(_17413__bF_buf7), .Y(_18085_) );
	OAI21X1 OAI21X1_3590 ( .gnd(gnd), .vdd(vdd), .A(_18084_), .B(_17412__bF_buf2), .C(_18085_), .Y(_18086_) );
	NOR2X1 NOR2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_18083_), .B(_18086_), .Y(_18087_) );
	INVX1 INVX1_2387 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_12_), .Y(_18088_) );
	NAND3X1 NAND3X1_3600 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(registers_r31_12_), .C(_17419__bF_buf2), .Y(_18089_) );
	OAI21X1 OAI21X1_3591 ( .gnd(gnd), .vdd(vdd), .A(_18088_), .B(_17418__bF_buf2), .C(_18089_), .Y(_18090_) );
	INVX1 INVX1_2388 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_12_), .Y(_18091_) );
	NAND3X1 NAND3X1_3601 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_12_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_18092_) );
	OAI21X1 OAI21X1_3592 ( .gnd(gnd), .vdd(vdd), .A(_18091_), .B(_17423__bF_buf2), .C(_18092_), .Y(_18093_) );
	NOR2X1 NOR2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_18090_), .B(_18093_), .Y(_18094_) );
	NAND2X1 NAND2X1_3438 ( .gnd(gnd), .vdd(vdd), .A(_18094_), .B(_18087_), .Y(_18095_) );
	NOR2X1 NOR2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_18095_), .B(_18080_), .Y(_18096_) );
	AOI22X1 AOI22X1_402 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf2), .B(registers_a2_12_), .C(registers_r1_12_), .D(_17431__bF_buf2), .Y(_18097_) );
	AOI22X1 AOI22X1_403 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf2), .B(registers_r4_12_), .C(registers_r5_12_), .D(_17436__bF_buf2), .Y(_18098_) );
	INVX1 INVX1_2389 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_12_), .Y(_18099_) );
	NAND3X1 NAND3X1_3602 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_12_), .B(_17432__bF_buf0), .C(_17392__bF_buf1), .Y(_18100_) );
	OAI21X1 OAI21X1_3593 ( .gnd(gnd), .vdd(vdd), .A(_18099_), .B(_17443__bF_buf2), .C(_18100_), .Y(_18101_) );
	AOI21X1 AOI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_12_), .B(_17440__bF_buf2), .C(_18101_), .Y(_18102_) );
	NAND3X1 NAND3X1_3603 ( .gnd(gnd), .vdd(vdd), .A(_18097_), .B(_18098_), .C(_18102_), .Y(_18103_) );
	INVX1 INVX1_2390 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_12_), .Y(_18104_) );
	INVX1 INVX1_2391 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_12_), .Y(_18105_) );
	OAI22X1 OAI22X1_252 ( .gnd(gnd), .vdd(vdd), .A(_18105_), .B(_17450__bF_buf2), .C(_18104_), .D(_17449__bF_buf2), .Y(_18106_) );
	INVX1 INVX1_2392 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_12_), .Y(_18107_) );
	INVX1 INVX1_2393 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_12_), .Y(_18108_) );
	OAI22X1 OAI22X1_253 ( .gnd(gnd), .vdd(vdd), .A(_18107_), .B(_17456__bF_buf2), .C(_18108_), .D(_17454__bF_buf2), .Y(_18109_) );
	NOR2X1 NOR2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_18109_), .B(_18106_), .Y(_18110_) );
	INVX1 INVX1_2394 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_12_), .Y(_18111_) );
	INVX1 INVX1_2395 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_12_), .Y(_18112_) );
	OAI22X1 OAI22X1_254 ( .gnd(gnd), .vdd(vdd), .A(_18111_), .B(_17461__bF_buf2), .C(_18112_), .D(_17462__bF_buf2), .Y(_18113_) );
	INVX1 INVX1_2396 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_12_), .Y(_18114_) );
	INVX1 INVX1_2397 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_12_), .Y(_18115_) );
	OAI22X1 OAI22X1_255 ( .gnd(gnd), .vdd(vdd), .A(_18115_), .B(_17467__bF_buf2), .C(_18114_), .D(_17466__bF_buf2), .Y(_18116_) );
	NOR2X1 NOR2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_18113_), .B(_18116_), .Y(_18117_) );
	NAND2X1 NAND2X1_3439 ( .gnd(gnd), .vdd(vdd), .A(_18110_), .B(_18117_), .Y(_18118_) );
	NOR2X1 NOR2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_18103_), .B(_18118_), .Y(_18119_) );
	NAND2X1 NAND2X1_3440 ( .gnd(gnd), .vdd(vdd), .A(_18119_), .B(_18096_), .Y(_428__12_) );
	NAND3X1 NAND3X1_3604 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_13_), .B(_17373__bF_buf4), .C(_17371__bF_buf4), .Y(_18120_) );
	NAND3X1 NAND3X1_3605 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_13_), .B(_17376__bF_buf4), .C(_17371__bF_buf3), .Y(_18121_) );
	NAND2X1 NAND2X1_3441 ( .gnd(gnd), .vdd(vdd), .A(_18120_), .B(_18121_), .Y(_18122_) );
	INVX1 INVX1_2398 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_13_), .Y(_18123_) );
	INVX1 INVX1_2399 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_13_), .Y(_18124_) );
	OAI22X1 OAI22X1_256 ( .gnd(gnd), .vdd(vdd), .A(_18123_), .B(_17384__bF_buf1), .C(_18124_), .D(_17383__bF_buf1), .Y(_18125_) );
	NOR2X1 NOR2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_18122_), .B(_18125_), .Y(_18126_) );
	INVX1 INVX1_2400 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_13_), .Y(_18127_) );
	INVX1 INVX1_2401 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_13_), .Y(_18128_) );
	OAI22X1 OAI22X1_257 ( .gnd(gnd), .vdd(vdd), .A(_18127_), .B(_17394__bF_buf1), .C(_18128_), .D(_17393__bF_buf1), .Y(_18129_) );
	INVX1 INVX1_2402 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_13_), .Y(_18130_) );
	INVX1 INVX1_2403 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_13_), .Y(_18131_) );
	OAI22X1 OAI22X1_258 ( .gnd(gnd), .vdd(vdd), .A(_18130_), .B(_17401__bF_buf1), .C(_18131_), .D(_17400__bF_buf1), .Y(_18132_) );
	NOR2X1 NOR2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_18132_), .B(_18129_), .Y(_18133_) );
	NAND2X1 NAND2X1_3442 ( .gnd(gnd), .vdd(vdd), .A(_18126_), .B(_18133_), .Y(_18134_) );
	INVX1 INVX1_2404 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_13_), .Y(_18135_) );
	INVX1 INVX1_2405 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_13_), .Y(_18136_) );
	OAI22X1 OAI22X1_259 ( .gnd(gnd), .vdd(vdd), .A(_18136_), .B(_17408__bF_buf1), .C(_18135_), .D(_17407__bF_buf1), .Y(_18137_) );
	INVX1 INVX1_2406 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_13_), .Y(_18138_) );
	NAND3X1 NAND3X1_3606 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_13_), .B(_17411__bF_buf0), .C(_17413__bF_buf5), .Y(_18139_) );
	OAI21X1 OAI21X1_3594 ( .gnd(gnd), .vdd(vdd), .A(_18138_), .B(_17412__bF_buf1), .C(_18139_), .Y(_18140_) );
	NOR2X1 NOR2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_18137_), .B(_18140_), .Y(_18141_) );
	INVX1 INVX1_2407 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_13_), .Y(_18142_) );
	NAND3X1 NAND3X1_3607 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(registers_r31_13_), .C(_17419__bF_buf1), .Y(_18143_) );
	OAI21X1 OAI21X1_3595 ( .gnd(gnd), .vdd(vdd), .A(_18142_), .B(_17418__bF_buf1), .C(_18143_), .Y(_18144_) );
	INVX1 INVX1_2408 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_13_), .Y(_18145_) );
	NAND3X1 NAND3X1_3608 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_13_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_18146_) );
	OAI21X1 OAI21X1_3596 ( .gnd(gnd), .vdd(vdd), .A(_18145_), .B(_17423__bF_buf1), .C(_18146_), .Y(_18147_) );
	NOR2X1 NOR2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_18144_), .B(_18147_), .Y(_18148_) );
	NAND2X1 NAND2X1_3443 ( .gnd(gnd), .vdd(vdd), .A(_18148_), .B(_18141_), .Y(_18149_) );
	NOR2X1 NOR2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_18149_), .B(_18134_), .Y(_18150_) );
	AOI22X1 AOI22X1_404 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf1), .B(registers_a2_13_), .C(registers_r1_13_), .D(_17431__bF_buf1), .Y(_18151_) );
	AOI22X1 AOI22X1_405 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf1), .B(registers_r4_13_), .C(registers_r5_13_), .D(_17436__bF_buf1), .Y(_18152_) );
	INVX1 INVX1_2409 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_13_), .Y(_18153_) );
	NAND3X1 NAND3X1_3609 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_13_), .B(_17432__bF_buf4), .C(_17392__bF_buf7), .Y(_18154_) );
	OAI21X1 OAI21X1_3597 ( .gnd(gnd), .vdd(vdd), .A(_18153_), .B(_17443__bF_buf1), .C(_18154_), .Y(_18155_) );
	AOI21X1 AOI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_13_), .B(_17440__bF_buf1), .C(_18155_), .Y(_18156_) );
	NAND3X1 NAND3X1_3610 ( .gnd(gnd), .vdd(vdd), .A(_18151_), .B(_18152_), .C(_18156_), .Y(_18157_) );
	INVX1 INVX1_2410 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_13_), .Y(_18158_) );
	INVX1 INVX1_2411 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_13_), .Y(_18159_) );
	OAI22X1 OAI22X1_260 ( .gnd(gnd), .vdd(vdd), .A(_18159_), .B(_17450__bF_buf1), .C(_18158_), .D(_17449__bF_buf1), .Y(_18160_) );
	INVX1 INVX1_2412 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_13_), .Y(_18161_) );
	INVX1 INVX1_2413 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_13_), .Y(_18162_) );
	OAI22X1 OAI22X1_261 ( .gnd(gnd), .vdd(vdd), .A(_18161_), .B(_17456__bF_buf1), .C(_18162_), .D(_17454__bF_buf1), .Y(_18163_) );
	NOR2X1 NOR2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_18163_), .B(_18160_), .Y(_18164_) );
	INVX1 INVX1_2414 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_13_), .Y(_18165_) );
	INVX1 INVX1_2415 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_13_), .Y(_18166_) );
	OAI22X1 OAI22X1_262 ( .gnd(gnd), .vdd(vdd), .A(_18165_), .B(_17461__bF_buf1), .C(_18166_), .D(_17462__bF_buf1), .Y(_18167_) );
	INVX1 INVX1_2416 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_13_), .Y(_18168_) );
	INVX1 INVX1_2417 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_13_), .Y(_18169_) );
	OAI22X1 OAI22X1_263 ( .gnd(gnd), .vdd(vdd), .A(_18169_), .B(_17467__bF_buf1), .C(_18168_), .D(_17466__bF_buf1), .Y(_18170_) );
	NOR2X1 NOR2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_18167_), .B(_18170_), .Y(_18171_) );
	NAND2X1 NAND2X1_3444 ( .gnd(gnd), .vdd(vdd), .A(_18164_), .B(_18171_), .Y(_18172_) );
	NOR2X1 NOR2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_18157_), .B(_18172_), .Y(_18173_) );
	NAND2X1 NAND2X1_3445 ( .gnd(gnd), .vdd(vdd), .A(_18173_), .B(_18150_), .Y(_428__13_) );
	NAND3X1 NAND3X1_3611 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_14_), .B(_17373__bF_buf3), .C(_17371__bF_buf2), .Y(_18174_) );
	NAND3X1 NAND3X1_3612 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_14_), .B(_17376__bF_buf3), .C(_17371__bF_buf1), .Y(_18175_) );
	NAND2X1 NAND2X1_3446 ( .gnd(gnd), .vdd(vdd), .A(_18174_), .B(_18175_), .Y(_18176_) );
	INVX1 INVX1_2418 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_14_), .Y(_18177_) );
	INVX1 INVX1_2419 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_14_), .Y(_18178_) );
	OAI22X1 OAI22X1_264 ( .gnd(gnd), .vdd(vdd), .A(_18177_), .B(_17384__bF_buf0), .C(_18178_), .D(_17383__bF_buf0), .Y(_18179_) );
	NOR2X1 NOR2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_18176_), .B(_18179_), .Y(_18180_) );
	INVX1 INVX1_2420 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_14_), .Y(_18181_) );
	INVX1 INVX1_2421 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_14_), .Y(_18182_) );
	OAI22X1 OAI22X1_265 ( .gnd(gnd), .vdd(vdd), .A(_18181_), .B(_17394__bF_buf0), .C(_18182_), .D(_17393__bF_buf0), .Y(_18183_) );
	INVX1 INVX1_2422 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_14_), .Y(_18184_) );
	INVX1 INVX1_2423 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_14_), .Y(_18185_) );
	OAI22X1 OAI22X1_266 ( .gnd(gnd), .vdd(vdd), .A(_18184_), .B(_17401__bF_buf0), .C(_18185_), .D(_17400__bF_buf0), .Y(_18186_) );
	NOR2X1 NOR2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_18186_), .B(_18183_), .Y(_18187_) );
	NAND2X1 NAND2X1_3447 ( .gnd(gnd), .vdd(vdd), .A(_18180_), .B(_18187_), .Y(_18188_) );
	INVX1 INVX1_2424 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_14_), .Y(_18189_) );
	INVX1 INVX1_2425 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_14_), .Y(_18190_) );
	OAI22X1 OAI22X1_267 ( .gnd(gnd), .vdd(vdd), .A(_18190_), .B(_17408__bF_buf0), .C(_18189_), .D(_17407__bF_buf0), .Y(_18191_) );
	INVX1 INVX1_2426 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_14_), .Y(_18192_) );
	NAND3X1 NAND3X1_3613 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_14_), .B(_17411__bF_buf5), .C(_17413__bF_buf3), .Y(_18193_) );
	OAI21X1 OAI21X1_3598 ( .gnd(gnd), .vdd(vdd), .A(_18192_), .B(_17412__bF_buf0), .C(_18193_), .Y(_18194_) );
	NOR2X1 NOR2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_18191_), .B(_18194_), .Y(_18195_) );
	INVX1 INVX1_2427 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_14_), .Y(_18196_) );
	NAND3X1 NAND3X1_3614 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(registers_r31_14_), .C(_17419__bF_buf0), .Y(_18197_) );
	OAI21X1 OAI21X1_3599 ( .gnd(gnd), .vdd(vdd), .A(_18196_), .B(_17418__bF_buf0), .C(_18197_), .Y(_18198_) );
	INVX1 INVX1_2428 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_14_), .Y(_18199_) );
	NAND3X1 NAND3X1_3615 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_14_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_18200_) );
	OAI21X1 OAI21X1_3600 ( .gnd(gnd), .vdd(vdd), .A(_18199_), .B(_17423__bF_buf0), .C(_18200_), .Y(_18201_) );
	NOR2X1 NOR2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_18198_), .B(_18201_), .Y(_18202_) );
	NAND2X1 NAND2X1_3448 ( .gnd(gnd), .vdd(vdd), .A(_18202_), .B(_18195_), .Y(_18203_) );
	NOR2X1 NOR2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_18203_), .B(_18188_), .Y(_18204_) );
	AOI22X1 AOI22X1_406 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf0), .B(registers_a2_14_), .C(registers_r1_14_), .D(_17431__bF_buf0), .Y(_18205_) );
	AOI22X1 AOI22X1_407 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf0), .B(registers_r4_14_), .C(registers_r5_14_), .D(_17436__bF_buf0), .Y(_18206_) );
	INVX1 INVX1_2429 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_14_), .Y(_18207_) );
	NAND3X1 NAND3X1_3616 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_14_), .B(_17432__bF_buf3), .C(_17392__bF_buf5), .Y(_18208_) );
	OAI21X1 OAI21X1_3601 ( .gnd(gnd), .vdd(vdd), .A(_18207_), .B(_17443__bF_buf0), .C(_18208_), .Y(_18209_) );
	AOI21X1 AOI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_14_), .B(_17440__bF_buf0), .C(_18209_), .Y(_18210_) );
	NAND3X1 NAND3X1_3617 ( .gnd(gnd), .vdd(vdd), .A(_18205_), .B(_18206_), .C(_18210_), .Y(_18211_) );
	INVX1 INVX1_2430 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_14_), .Y(_18212_) );
	INVX1 INVX1_2431 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_14_), .Y(_18213_) );
	OAI22X1 OAI22X1_268 ( .gnd(gnd), .vdd(vdd), .A(_18213_), .B(_17450__bF_buf0), .C(_18212_), .D(_17449__bF_buf0), .Y(_18214_) );
	INVX1 INVX1_2432 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_14_), .Y(_18215_) );
	INVX1 INVX1_2433 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_14_), .Y(_18216_) );
	OAI22X1 OAI22X1_269 ( .gnd(gnd), .vdd(vdd), .A(_18215_), .B(_17456__bF_buf0), .C(_18216_), .D(_17454__bF_buf0), .Y(_18217_) );
	NOR2X1 NOR2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_18217_), .B(_18214_), .Y(_18218_) );
	INVX1 INVX1_2434 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_14_), .Y(_18219_) );
	INVX1 INVX1_2435 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_14_), .Y(_18220_) );
	OAI22X1 OAI22X1_270 ( .gnd(gnd), .vdd(vdd), .A(_18219_), .B(_17461__bF_buf0), .C(_18220_), .D(_17462__bF_buf0), .Y(_18221_) );
	INVX1 INVX1_2436 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_14_), .Y(_18222_) );
	INVX1 INVX1_2437 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_14_), .Y(_18223_) );
	OAI22X1 OAI22X1_271 ( .gnd(gnd), .vdd(vdd), .A(_18223_), .B(_17467__bF_buf0), .C(_18222_), .D(_17466__bF_buf0), .Y(_18224_) );
	NOR2X1 NOR2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_18221_), .B(_18224_), .Y(_18225_) );
	NAND2X1 NAND2X1_3449 ( .gnd(gnd), .vdd(vdd), .A(_18218_), .B(_18225_), .Y(_18226_) );
	NOR2X1 NOR2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_18211_), .B(_18226_), .Y(_18227_) );
	NAND2X1 NAND2X1_3450 ( .gnd(gnd), .vdd(vdd), .A(_18227_), .B(_18204_), .Y(_428__14_) );
	NAND3X1 NAND3X1_3618 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_15_), .B(_17373__bF_buf2), .C(_17371__bF_buf0), .Y(_18228_) );
	NAND3X1 NAND3X1_3619 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_15_), .B(_17376__bF_buf2), .C(_17371__bF_buf7), .Y(_18229_) );
	NAND2X1 NAND2X1_3451 ( .gnd(gnd), .vdd(vdd), .A(_18228_), .B(_18229_), .Y(_18230_) );
	INVX1 INVX1_2438 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_15_), .Y(_18231_) );
	INVX1 INVX1_2439 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_15_), .Y(_18232_) );
	OAI22X1 OAI22X1_272 ( .gnd(gnd), .vdd(vdd), .A(_18231_), .B(_17384__bF_buf4), .C(_18232_), .D(_17383__bF_buf4), .Y(_18233_) );
	NOR2X1 NOR2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_18230_), .B(_18233_), .Y(_18234_) );
	INVX1 INVX1_2440 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_15_), .Y(_18235_) );
	INVX1 INVX1_2441 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_15_), .Y(_18236_) );
	OAI22X1 OAI22X1_273 ( .gnd(gnd), .vdd(vdd), .A(_18235_), .B(_17394__bF_buf4), .C(_18236_), .D(_17393__bF_buf4), .Y(_18237_) );
	INVX1 INVX1_2442 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_15_), .Y(_18238_) );
	INVX1 INVX1_2443 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_15_), .Y(_18239_) );
	OAI22X1 OAI22X1_274 ( .gnd(gnd), .vdd(vdd), .A(_18238_), .B(_17401__bF_buf4), .C(_18239_), .D(_17400__bF_buf4), .Y(_18240_) );
	NOR2X1 NOR2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_18240_), .B(_18237_), .Y(_18241_) );
	NAND2X1 NAND2X1_3452 ( .gnd(gnd), .vdd(vdd), .A(_18234_), .B(_18241_), .Y(_18242_) );
	INVX1 INVX1_2444 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_15_), .Y(_18243_) );
	INVX1 INVX1_2445 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_15_), .Y(_18244_) );
	OAI22X1 OAI22X1_275 ( .gnd(gnd), .vdd(vdd), .A(_18244_), .B(_17408__bF_buf4), .C(_18243_), .D(_17407__bF_buf4), .Y(_18245_) );
	INVX1 INVX1_2446 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_15_), .Y(_18246_) );
	NAND3X1 NAND3X1_3620 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_15_), .B(_17411__bF_buf4), .C(_17413__bF_buf1), .Y(_18247_) );
	OAI21X1 OAI21X1_3602 ( .gnd(gnd), .vdd(vdd), .A(_18246_), .B(_17412__bF_buf4), .C(_18247_), .Y(_18248_) );
	NOR2X1 NOR2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_18245_), .B(_18248_), .Y(_18249_) );
	INVX1 INVX1_2447 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_15_), .Y(_18250_) );
	NAND3X1 NAND3X1_3621 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(registers_r31_15_), .C(_17419__bF_buf4), .Y(_18251_) );
	OAI21X1 OAI21X1_3603 ( .gnd(gnd), .vdd(vdd), .A(_18250_), .B(_17418__bF_buf4), .C(_18251_), .Y(_18252_) );
	INVX1 INVX1_2448 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_15_), .Y(_18253_) );
	NAND3X1 NAND3X1_3622 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_15_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_18254_) );
	OAI21X1 OAI21X1_3604 ( .gnd(gnd), .vdd(vdd), .A(_18253_), .B(_17423__bF_buf4), .C(_18254_), .Y(_18255_) );
	NOR2X1 NOR2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_18252_), .B(_18255_), .Y(_18256_) );
	NAND2X1 NAND2X1_3453 ( .gnd(gnd), .vdd(vdd), .A(_18256_), .B(_18249_), .Y(_18257_) );
	NOR2X1 NOR2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_18257_), .B(_18242_), .Y(_18258_) );
	AOI22X1 AOI22X1_408 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_15_), .C(registers_r1_15_), .D(_17431__bF_buf4), .Y(_18259_) );
	AOI22X1 AOI22X1_409 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_15_), .C(registers_r5_15_), .D(_17436__bF_buf4), .Y(_18260_) );
	INVX1 INVX1_2449 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_15_), .Y(_18261_) );
	NAND3X1 NAND3X1_3623 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_15_), .B(_17432__bF_buf2), .C(_17392__bF_buf3), .Y(_18262_) );
	OAI21X1 OAI21X1_3605 ( .gnd(gnd), .vdd(vdd), .A(_18261_), .B(_17443__bF_buf4), .C(_18262_), .Y(_18263_) );
	AOI21X1 AOI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_15_), .B(_17440__bF_buf4), .C(_18263_), .Y(_18264_) );
	NAND3X1 NAND3X1_3624 ( .gnd(gnd), .vdd(vdd), .A(_18259_), .B(_18260_), .C(_18264_), .Y(_18265_) );
	INVX1 INVX1_2450 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_15_), .Y(_18266_) );
	INVX1 INVX1_2451 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_15_), .Y(_18267_) );
	OAI22X1 OAI22X1_276 ( .gnd(gnd), .vdd(vdd), .A(_18267_), .B(_17450__bF_buf4), .C(_18266_), .D(_17449__bF_buf4), .Y(_18268_) );
	INVX1 INVX1_2452 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_15_), .Y(_18269_) );
	INVX1 INVX1_2453 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_15_), .Y(_18270_) );
	OAI22X1 OAI22X1_277 ( .gnd(gnd), .vdd(vdd), .A(_18269_), .B(_17456__bF_buf4), .C(_18270_), .D(_17454__bF_buf4), .Y(_18271_) );
	NOR2X1 NOR2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_18271_), .B(_18268_), .Y(_18272_) );
	INVX1 INVX1_2454 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_15_), .Y(_18273_) );
	INVX1 INVX1_2455 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_15_), .Y(_18274_) );
	OAI22X1 OAI22X1_278 ( .gnd(gnd), .vdd(vdd), .A(_18273_), .B(_17461__bF_buf4), .C(_18274_), .D(_17462__bF_buf4), .Y(_18275_) );
	INVX1 INVX1_2456 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_15_), .Y(_18276_) );
	INVX1 INVX1_2457 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_15_), .Y(_18277_) );
	OAI22X1 OAI22X1_279 ( .gnd(gnd), .vdd(vdd), .A(_18277_), .B(_17467__bF_buf4), .C(_18276_), .D(_17466__bF_buf4), .Y(_18278_) );
	NOR2X1 NOR2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_18275_), .B(_18278_), .Y(_18279_) );
	NAND2X1 NAND2X1_3454 ( .gnd(gnd), .vdd(vdd), .A(_18272_), .B(_18279_), .Y(_18280_) );
	NOR2X1 NOR2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_18265_), .B(_18280_), .Y(_18281_) );
	NAND2X1 NAND2X1_3455 ( .gnd(gnd), .vdd(vdd), .A(_18281_), .B(_18258_), .Y(_428__15_) );
	NAND3X1 NAND3X1_3625 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_16_), .B(_17373__bF_buf1), .C(_17371__bF_buf6), .Y(_18282_) );
	NAND3X1 NAND3X1_3626 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_16_), .B(_17376__bF_buf1), .C(_17371__bF_buf5), .Y(_18283_) );
	NAND2X1 NAND2X1_3456 ( .gnd(gnd), .vdd(vdd), .A(_18282_), .B(_18283_), .Y(_18284_) );
	INVX1 INVX1_2458 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_16_), .Y(_18285_) );
	INVX1 INVX1_2459 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_16_), .Y(_18286_) );
	OAI22X1 OAI22X1_280 ( .gnd(gnd), .vdd(vdd), .A(_18285_), .B(_17384__bF_buf3), .C(_18286_), .D(_17383__bF_buf3), .Y(_18287_) );
	NOR2X1 NOR2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_18284_), .B(_18287_), .Y(_18288_) );
	INVX1 INVX1_2460 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_16_), .Y(_18289_) );
	INVX1 INVX1_2461 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_16_), .Y(_18290_) );
	OAI22X1 OAI22X1_281 ( .gnd(gnd), .vdd(vdd), .A(_18289_), .B(_17394__bF_buf3), .C(_18290_), .D(_17393__bF_buf3), .Y(_18291_) );
	INVX1 INVX1_2462 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_16_), .Y(_18292_) );
	INVX1 INVX1_2463 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_16_), .Y(_18293_) );
	OAI22X1 OAI22X1_282 ( .gnd(gnd), .vdd(vdd), .A(_18292_), .B(_17401__bF_buf3), .C(_18293_), .D(_17400__bF_buf3), .Y(_18294_) );
	NOR2X1 NOR2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_18294_), .B(_18291_), .Y(_18295_) );
	NAND2X1 NAND2X1_3457 ( .gnd(gnd), .vdd(vdd), .A(_18288_), .B(_18295_), .Y(_18296_) );
	INVX1 INVX1_2464 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_16_), .Y(_18297_) );
	INVX1 INVX1_2465 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_16_), .Y(_18298_) );
	OAI22X1 OAI22X1_283 ( .gnd(gnd), .vdd(vdd), .A(_18298_), .B(_17408__bF_buf3), .C(_18297_), .D(_17407__bF_buf3), .Y(_18299_) );
	INVX1 INVX1_2466 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_16_), .Y(_18300_) );
	NAND3X1 NAND3X1_3627 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_16_), .B(_17411__bF_buf3), .C(_17413__bF_buf7), .Y(_18301_) );
	OAI21X1 OAI21X1_3606 ( .gnd(gnd), .vdd(vdd), .A(_18300_), .B(_17412__bF_buf3), .C(_18301_), .Y(_18302_) );
	NOR2X1 NOR2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_18299_), .B(_18302_), .Y(_18303_) );
	INVX1 INVX1_2467 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_16_), .Y(_18304_) );
	NAND3X1 NAND3X1_3628 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(registers_r31_16_), .C(_17419__bF_buf3), .Y(_18305_) );
	OAI21X1 OAI21X1_3607 ( .gnd(gnd), .vdd(vdd), .A(_18304_), .B(_17418__bF_buf3), .C(_18305_), .Y(_18306_) );
	INVX1 INVX1_2468 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_16_), .Y(_18307_) );
	NAND3X1 NAND3X1_3629 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_16_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_18308_) );
	OAI21X1 OAI21X1_3608 ( .gnd(gnd), .vdd(vdd), .A(_18307_), .B(_17423__bF_buf3), .C(_18308_), .Y(_18309_) );
	NOR2X1 NOR2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_18306_), .B(_18309_), .Y(_18310_) );
	NAND2X1 NAND2X1_3458 ( .gnd(gnd), .vdd(vdd), .A(_18310_), .B(_18303_), .Y(_18311_) );
	NOR2X1 NOR2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_18311_), .B(_18296_), .Y(_18312_) );
	AOI22X1 AOI22X1_410 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_16_), .C(registers_r1_16_), .D(_17431__bF_buf3), .Y(_18313_) );
	AOI22X1 AOI22X1_411 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_16_), .C(registers_r5_16_), .D(_17436__bF_buf3), .Y(_18314_) );
	INVX1 INVX1_2469 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_16_), .Y(_18315_) );
	NAND3X1 NAND3X1_3630 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_16_), .B(_17432__bF_buf1), .C(_17392__bF_buf1), .Y(_18316_) );
	OAI21X1 OAI21X1_3609 ( .gnd(gnd), .vdd(vdd), .A(_18315_), .B(_17443__bF_buf3), .C(_18316_), .Y(_18317_) );
	AOI21X1 AOI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_16_), .B(_17440__bF_buf3), .C(_18317_), .Y(_18318_) );
	NAND3X1 NAND3X1_3631 ( .gnd(gnd), .vdd(vdd), .A(_18313_), .B(_18314_), .C(_18318_), .Y(_18319_) );
	INVX1 INVX1_2470 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_16_), .Y(_18320_) );
	INVX1 INVX1_2471 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_16_), .Y(_18321_) );
	OAI22X1 OAI22X1_284 ( .gnd(gnd), .vdd(vdd), .A(_18321_), .B(_17450__bF_buf3), .C(_18320_), .D(_17449__bF_buf3), .Y(_18322_) );
	INVX1 INVX1_2472 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_16_), .Y(_18323_) );
	INVX1 INVX1_2473 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_16_), .Y(_18324_) );
	OAI22X1 OAI22X1_285 ( .gnd(gnd), .vdd(vdd), .A(_18323_), .B(_17456__bF_buf3), .C(_18324_), .D(_17454__bF_buf3), .Y(_18325_) );
	NOR2X1 NOR2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_18325_), .B(_18322_), .Y(_18326_) );
	INVX1 INVX1_2474 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_16_), .Y(_18327_) );
	INVX1 INVX1_2475 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_16_), .Y(_18328_) );
	OAI22X1 OAI22X1_286 ( .gnd(gnd), .vdd(vdd), .A(_18327_), .B(_17461__bF_buf3), .C(_18328_), .D(_17462__bF_buf3), .Y(_18329_) );
	INVX1 INVX1_2476 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_16_), .Y(_18330_) );
	INVX1 INVX1_2477 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_16_), .Y(_18331_) );
	OAI22X1 OAI22X1_287 ( .gnd(gnd), .vdd(vdd), .A(_18331_), .B(_17467__bF_buf3), .C(_18330_), .D(_17466__bF_buf3), .Y(_18332_) );
	NOR2X1 NOR2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_18329_), .B(_18332_), .Y(_18333_) );
	NAND2X1 NAND2X1_3459 ( .gnd(gnd), .vdd(vdd), .A(_18326_), .B(_18333_), .Y(_18334_) );
	NOR2X1 NOR2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_18319_), .B(_18334_), .Y(_18335_) );
	NAND2X1 NAND2X1_3460 ( .gnd(gnd), .vdd(vdd), .A(_18335_), .B(_18312_), .Y(_428__16_) );
	NAND3X1 NAND3X1_3632 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_17_), .B(_17373__bF_buf0), .C(_17371__bF_buf4), .Y(_18336_) );
	NAND3X1 NAND3X1_3633 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_17_), .B(_17376__bF_buf0), .C(_17371__bF_buf3), .Y(_18337_) );
	NAND2X1 NAND2X1_3461 ( .gnd(gnd), .vdd(vdd), .A(_18336_), .B(_18337_), .Y(_18338_) );
	INVX1 INVX1_2478 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_17_), .Y(_18339_) );
	INVX1 INVX1_2479 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_17_), .Y(_18340_) );
	OAI22X1 OAI22X1_288 ( .gnd(gnd), .vdd(vdd), .A(_18339_), .B(_17384__bF_buf2), .C(_18340_), .D(_17383__bF_buf2), .Y(_18341_) );
	NOR2X1 NOR2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_18338_), .B(_18341_), .Y(_18342_) );
	INVX1 INVX1_2480 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_17_), .Y(_18343_) );
	INVX1 INVX1_2481 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_17_), .Y(_18344_) );
	OAI22X1 OAI22X1_289 ( .gnd(gnd), .vdd(vdd), .A(_18343_), .B(_17394__bF_buf2), .C(_18344_), .D(_17393__bF_buf2), .Y(_18345_) );
	INVX1 INVX1_2482 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_17_), .Y(_18346_) );
	INVX1 INVX1_2483 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_17_), .Y(_18347_) );
	OAI22X1 OAI22X1_290 ( .gnd(gnd), .vdd(vdd), .A(_18346_), .B(_17401__bF_buf2), .C(_18347_), .D(_17400__bF_buf2), .Y(_18348_) );
	NOR2X1 NOR2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_18348_), .B(_18345_), .Y(_18349_) );
	NAND2X1 NAND2X1_3462 ( .gnd(gnd), .vdd(vdd), .A(_18342_), .B(_18349_), .Y(_18350_) );
	INVX1 INVX1_2484 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_17_), .Y(_18351_) );
	INVX1 INVX1_2485 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_17_), .Y(_18352_) );
	OAI22X1 OAI22X1_291 ( .gnd(gnd), .vdd(vdd), .A(_18352_), .B(_17408__bF_buf2), .C(_18351_), .D(_17407__bF_buf2), .Y(_18353_) );
	INVX1 INVX1_2486 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_17_), .Y(_18354_) );
	NAND3X1 NAND3X1_3634 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_17_), .B(_17411__bF_buf2), .C(_17413__bF_buf5), .Y(_18355_) );
	OAI21X1 OAI21X1_3610 ( .gnd(gnd), .vdd(vdd), .A(_18354_), .B(_17412__bF_buf2), .C(_18355_), .Y(_18356_) );
	NOR2X1 NOR2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_18353_), .B(_18356_), .Y(_18357_) );
	INVX1 INVX1_2487 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_17_), .Y(_18358_) );
	NAND3X1 NAND3X1_3635 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(registers_r31_17_), .C(_17419__bF_buf2), .Y(_18359_) );
	OAI21X1 OAI21X1_3611 ( .gnd(gnd), .vdd(vdd), .A(_18358_), .B(_17418__bF_buf2), .C(_18359_), .Y(_18360_) );
	INVX1 INVX1_2488 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_17_), .Y(_18361_) );
	NAND3X1 NAND3X1_3636 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_17_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_18362_) );
	OAI21X1 OAI21X1_3612 ( .gnd(gnd), .vdd(vdd), .A(_18361_), .B(_17423__bF_buf2), .C(_18362_), .Y(_18363_) );
	NOR2X1 NOR2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_18360_), .B(_18363_), .Y(_18364_) );
	NAND2X1 NAND2X1_3463 ( .gnd(gnd), .vdd(vdd), .A(_18364_), .B(_18357_), .Y(_18365_) );
	NOR2X1 NOR2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_18365_), .B(_18350_), .Y(_18366_) );
	AOI22X1 AOI22X1_412 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf2), .B(registers_a2_17_), .C(registers_r1_17_), .D(_17431__bF_buf2), .Y(_18367_) );
	AOI22X1 AOI22X1_413 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf2), .B(registers_r4_17_), .C(registers_r5_17_), .D(_17436__bF_buf2), .Y(_18368_) );
	INVX1 INVX1_2489 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_17_), .Y(_18369_) );
	NAND3X1 NAND3X1_3637 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_17_), .B(_17432__bF_buf0), .C(_17392__bF_buf7), .Y(_18370_) );
	OAI21X1 OAI21X1_3613 ( .gnd(gnd), .vdd(vdd), .A(_18369_), .B(_17443__bF_buf2), .C(_18370_), .Y(_18371_) );
	AOI21X1 AOI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_17_), .B(_17440__bF_buf2), .C(_18371_), .Y(_18372_) );
	NAND3X1 NAND3X1_3638 ( .gnd(gnd), .vdd(vdd), .A(_18367_), .B(_18368_), .C(_18372_), .Y(_18373_) );
	INVX1 INVX1_2490 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_17_), .Y(_18374_) );
	INVX1 INVX1_2491 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_17_), .Y(_18375_) );
	OAI22X1 OAI22X1_292 ( .gnd(gnd), .vdd(vdd), .A(_18375_), .B(_17450__bF_buf2), .C(_18374_), .D(_17449__bF_buf2), .Y(_18376_) );
	INVX1 INVX1_2492 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_17_), .Y(_18377_) );
	INVX1 INVX1_2493 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_17_), .Y(_18378_) );
	OAI22X1 OAI22X1_293 ( .gnd(gnd), .vdd(vdd), .A(_18377_), .B(_17456__bF_buf2), .C(_18378_), .D(_17454__bF_buf2), .Y(_18379_) );
	NOR2X1 NOR2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_18379_), .B(_18376_), .Y(_18380_) );
	INVX1 INVX1_2494 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_17_), .Y(_18381_) );
	INVX1 INVX1_2495 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_17_), .Y(_18382_) );
	OAI22X1 OAI22X1_294 ( .gnd(gnd), .vdd(vdd), .A(_18381_), .B(_17461__bF_buf2), .C(_18382_), .D(_17462__bF_buf2), .Y(_18383_) );
	INVX1 INVX1_2496 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_17_), .Y(_18384_) );
	INVX1 INVX1_2497 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_17_), .Y(_18385_) );
	OAI22X1 OAI22X1_295 ( .gnd(gnd), .vdd(vdd), .A(_18385_), .B(_17467__bF_buf2), .C(_18384_), .D(_17466__bF_buf2), .Y(_18386_) );
	NOR2X1 NOR2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_18383_), .B(_18386_), .Y(_18387_) );
	NAND2X1 NAND2X1_3464 ( .gnd(gnd), .vdd(vdd), .A(_18380_), .B(_18387_), .Y(_18388_) );
	NOR2X1 NOR2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_18373_), .B(_18388_), .Y(_18389_) );
	NAND2X1 NAND2X1_3465 ( .gnd(gnd), .vdd(vdd), .A(_18389_), .B(_18366_), .Y(_428__17_) );
	NAND3X1 NAND3X1_3639 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_18_), .B(_17373__bF_buf5), .C(_17371__bF_buf2), .Y(_18390_) );
	NAND3X1 NAND3X1_3640 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_18_), .B(_17376__bF_buf5), .C(_17371__bF_buf1), .Y(_18391_) );
	NAND2X1 NAND2X1_3466 ( .gnd(gnd), .vdd(vdd), .A(_18390_), .B(_18391_), .Y(_18392_) );
	INVX1 INVX1_2498 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_18_), .Y(_18393_) );
	INVX1 INVX1_2499 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_18_), .Y(_18394_) );
	OAI22X1 OAI22X1_296 ( .gnd(gnd), .vdd(vdd), .A(_18393_), .B(_17384__bF_buf1), .C(_18394_), .D(_17383__bF_buf1), .Y(_18395_) );
	NOR2X1 NOR2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_18392_), .B(_18395_), .Y(_18396_) );
	INVX1 INVX1_2500 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_18_), .Y(_18397_) );
	INVX1 INVX1_2501 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_18_), .Y(_18398_) );
	OAI22X1 OAI22X1_297 ( .gnd(gnd), .vdd(vdd), .A(_18397_), .B(_17394__bF_buf1), .C(_18398_), .D(_17393__bF_buf1), .Y(_18399_) );
	INVX1 INVX1_2502 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_18_), .Y(_18400_) );
	INVX1 INVX1_2503 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_18_), .Y(_18401_) );
	OAI22X1 OAI22X1_298 ( .gnd(gnd), .vdd(vdd), .A(_18400_), .B(_17401__bF_buf1), .C(_18401_), .D(_17400__bF_buf1), .Y(_18402_) );
	NOR2X1 NOR2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_18402_), .B(_18399_), .Y(_18403_) );
	NAND2X1 NAND2X1_3467 ( .gnd(gnd), .vdd(vdd), .A(_18396_), .B(_18403_), .Y(_18404_) );
	INVX1 INVX1_2504 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_18_), .Y(_18405_) );
	INVX1 INVX1_2505 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_18_), .Y(_18406_) );
	OAI22X1 OAI22X1_299 ( .gnd(gnd), .vdd(vdd), .A(_18406_), .B(_17408__bF_buf1), .C(_18405_), .D(_17407__bF_buf1), .Y(_18407_) );
	INVX1 INVX1_2506 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_18_), .Y(_18408_) );
	NAND3X1 NAND3X1_3641 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_18_), .B(_17411__bF_buf1), .C(_17413__bF_buf3), .Y(_18409_) );
	OAI21X1 OAI21X1_3614 ( .gnd(gnd), .vdd(vdd), .A(_18408_), .B(_17412__bF_buf1), .C(_18409_), .Y(_18410_) );
	NOR2X1 NOR2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_18407_), .B(_18410_), .Y(_18411_) );
	INVX1 INVX1_2507 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_18_), .Y(_18412_) );
	NAND3X1 NAND3X1_3642 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .B(registers_r31_18_), .C(_17419__bF_buf1), .Y(_18413_) );
	OAI21X1 OAI21X1_3615 ( .gnd(gnd), .vdd(vdd), .A(_18412_), .B(_17418__bF_buf1), .C(_18413_), .Y(_18414_) );
	INVX1 INVX1_2508 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_18_), .Y(_18415_) );
	NAND3X1 NAND3X1_3643 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_18_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_18416_) );
	OAI21X1 OAI21X1_3616 ( .gnd(gnd), .vdd(vdd), .A(_18415_), .B(_17423__bF_buf1), .C(_18416_), .Y(_18417_) );
	NOR2X1 NOR2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_18414_), .B(_18417_), .Y(_18418_) );
	NAND2X1 NAND2X1_3468 ( .gnd(gnd), .vdd(vdd), .A(_18418_), .B(_18411_), .Y(_18419_) );
	NOR2X1 NOR2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_18419_), .B(_18404_), .Y(_18420_) );
	AOI22X1 AOI22X1_414 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf1), .B(registers_a2_18_), .C(registers_r1_18_), .D(_17431__bF_buf1), .Y(_18421_) );
	AOI22X1 AOI22X1_415 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf1), .B(registers_r4_18_), .C(registers_r5_18_), .D(_17436__bF_buf1), .Y(_18422_) );
	INVX1 INVX1_2509 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_18_), .Y(_18423_) );
	NAND3X1 NAND3X1_3644 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_18_), .B(_17432__bF_buf4), .C(_17392__bF_buf5), .Y(_18424_) );
	OAI21X1 OAI21X1_3617 ( .gnd(gnd), .vdd(vdd), .A(_18423_), .B(_17443__bF_buf1), .C(_18424_), .Y(_18425_) );
	AOI21X1 AOI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_18_), .B(_17440__bF_buf1), .C(_18425_), .Y(_18426_) );
	NAND3X1 NAND3X1_3645 ( .gnd(gnd), .vdd(vdd), .A(_18421_), .B(_18422_), .C(_18426_), .Y(_18427_) );
	INVX1 INVX1_2510 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_18_), .Y(_18428_) );
	INVX1 INVX1_2511 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_18_), .Y(_18429_) );
	OAI22X1 OAI22X1_300 ( .gnd(gnd), .vdd(vdd), .A(_18429_), .B(_17450__bF_buf1), .C(_18428_), .D(_17449__bF_buf1), .Y(_18430_) );
	INVX1 INVX1_2512 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_18_), .Y(_18431_) );
	INVX1 INVX1_2513 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_18_), .Y(_18432_) );
	OAI22X1 OAI22X1_301 ( .gnd(gnd), .vdd(vdd), .A(_18431_), .B(_17456__bF_buf1), .C(_18432_), .D(_17454__bF_buf1), .Y(_18433_) );
	NOR2X1 NOR2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_18433_), .B(_18430_), .Y(_18434_) );
	INVX1 INVX1_2514 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_18_), .Y(_18435_) );
	INVX1 INVX1_2515 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_18_), .Y(_18436_) );
	OAI22X1 OAI22X1_302 ( .gnd(gnd), .vdd(vdd), .A(_18435_), .B(_17461__bF_buf1), .C(_18436_), .D(_17462__bF_buf1), .Y(_18437_) );
	INVX1 INVX1_2516 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_18_), .Y(_18438_) );
	INVX1 INVX1_2517 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_18_), .Y(_18439_) );
	OAI22X1 OAI22X1_303 ( .gnd(gnd), .vdd(vdd), .A(_18439_), .B(_17467__bF_buf1), .C(_18438_), .D(_17466__bF_buf1), .Y(_18440_) );
	NOR2X1 NOR2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_18437_), .B(_18440_), .Y(_18441_) );
	NAND2X1 NAND2X1_3469 ( .gnd(gnd), .vdd(vdd), .A(_18434_), .B(_18441_), .Y(_18442_) );
	NOR2X1 NOR2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_18427_), .B(_18442_), .Y(_18443_) );
	NAND2X1 NAND2X1_3470 ( .gnd(gnd), .vdd(vdd), .A(_18443_), .B(_18420_), .Y(_428__18_) );
	NAND3X1 NAND3X1_3646 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_19_), .B(_17373__bF_buf4), .C(_17371__bF_buf0), .Y(_18444_) );
	NAND3X1 NAND3X1_3647 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_19_), .B(_17376__bF_buf4), .C(_17371__bF_buf7), .Y(_18445_) );
	NAND2X1 NAND2X1_3471 ( .gnd(gnd), .vdd(vdd), .A(_18444_), .B(_18445_), .Y(_18446_) );
	INVX1 INVX1_2518 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_19_), .Y(_18447_) );
	INVX1 INVX1_2519 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_19_), .Y(_18448_) );
	OAI22X1 OAI22X1_304 ( .gnd(gnd), .vdd(vdd), .A(_18447_), .B(_17384__bF_buf0), .C(_18448_), .D(_17383__bF_buf0), .Y(_18449_) );
	NOR2X1 NOR2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_18446_), .B(_18449_), .Y(_18450_) );
	INVX1 INVX1_2520 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_19_), .Y(_18451_) );
	INVX1 INVX1_2521 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_19_), .Y(_18452_) );
	OAI22X1 OAI22X1_305 ( .gnd(gnd), .vdd(vdd), .A(_18451_), .B(_17394__bF_buf0), .C(_18452_), .D(_17393__bF_buf0), .Y(_18453_) );
	INVX1 INVX1_2522 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_19_), .Y(_18454_) );
	INVX1 INVX1_2523 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_19_), .Y(_18455_) );
	OAI22X1 OAI22X1_306 ( .gnd(gnd), .vdd(vdd), .A(_18454_), .B(_17401__bF_buf0), .C(_18455_), .D(_17400__bF_buf0), .Y(_18456_) );
	NOR2X1 NOR2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_18456_), .B(_18453_), .Y(_18457_) );
	NAND2X1 NAND2X1_3472 ( .gnd(gnd), .vdd(vdd), .A(_18450_), .B(_18457_), .Y(_18458_) );
	INVX1 INVX1_2524 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_19_), .Y(_18459_) );
	INVX1 INVX1_2525 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_19_), .Y(_18460_) );
	OAI22X1 OAI22X1_307 ( .gnd(gnd), .vdd(vdd), .A(_18460_), .B(_17408__bF_buf0), .C(_18459_), .D(_17407__bF_buf0), .Y(_18461_) );
	INVX1 INVX1_2526 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_19_), .Y(_18462_) );
	NAND3X1 NAND3X1_3648 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_19_), .B(_17411__bF_buf0), .C(_17413__bF_buf1), .Y(_18463_) );
	OAI21X1 OAI21X1_3618 ( .gnd(gnd), .vdd(vdd), .A(_18462_), .B(_17412__bF_buf0), .C(_18463_), .Y(_18464_) );
	NOR2X1 NOR2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_18461_), .B(_18464_), .Y(_18465_) );
	INVX1 INVX1_2527 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_19_), .Y(_18466_) );
	NAND3X1 NAND3X1_3649 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(registers_r31_19_), .C(_17419__bF_buf0), .Y(_18467_) );
	OAI21X1 OAI21X1_3619 ( .gnd(gnd), .vdd(vdd), .A(_18466_), .B(_17418__bF_buf0), .C(_18467_), .Y(_18468_) );
	INVX1 INVX1_2528 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_19_), .Y(_18469_) );
	NAND3X1 NAND3X1_3650 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_19_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_18470_) );
	OAI21X1 OAI21X1_3620 ( .gnd(gnd), .vdd(vdd), .A(_18469_), .B(_17423__bF_buf0), .C(_18470_), .Y(_18471_) );
	NOR2X1 NOR2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_18468_), .B(_18471_), .Y(_18472_) );
	NAND2X1 NAND2X1_3473 ( .gnd(gnd), .vdd(vdd), .A(_18472_), .B(_18465_), .Y(_18473_) );
	NOR2X1 NOR2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_18473_), .B(_18458_), .Y(_18474_) );
	AOI22X1 AOI22X1_416 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf0), .B(registers_a2_19_), .C(registers_r1_19_), .D(_17431__bF_buf0), .Y(_18475_) );
	AOI22X1 AOI22X1_417 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf0), .B(registers_r4_19_), .C(registers_r5_19_), .D(_17436__bF_buf0), .Y(_18476_) );
	INVX1 INVX1_2529 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_19_), .Y(_18477_) );
	NAND3X1 NAND3X1_3651 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_19_), .B(_17432__bF_buf3), .C(_17392__bF_buf3), .Y(_18478_) );
	OAI21X1 OAI21X1_3621 ( .gnd(gnd), .vdd(vdd), .A(_18477_), .B(_17443__bF_buf0), .C(_18478_), .Y(_18479_) );
	AOI21X1 AOI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_19_), .B(_17440__bF_buf0), .C(_18479_), .Y(_18480_) );
	NAND3X1 NAND3X1_3652 ( .gnd(gnd), .vdd(vdd), .A(_18475_), .B(_18476_), .C(_18480_), .Y(_18481_) );
	INVX1 INVX1_2530 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_19_), .Y(_18482_) );
	INVX1 INVX1_2531 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_19_), .Y(_18483_) );
	OAI22X1 OAI22X1_308 ( .gnd(gnd), .vdd(vdd), .A(_18483_), .B(_17450__bF_buf0), .C(_18482_), .D(_17449__bF_buf0), .Y(_18484_) );
	INVX1 INVX1_2532 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_19_), .Y(_18485_) );
	INVX1 INVX1_2533 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_19_), .Y(_18486_) );
	OAI22X1 OAI22X1_309 ( .gnd(gnd), .vdd(vdd), .A(_18485_), .B(_17456__bF_buf0), .C(_18486_), .D(_17454__bF_buf0), .Y(_18487_) );
	NOR2X1 NOR2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_18487_), .B(_18484_), .Y(_18488_) );
	INVX1 INVX1_2534 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_19_), .Y(_18489_) );
	INVX1 INVX1_2535 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_19_), .Y(_18490_) );
	OAI22X1 OAI22X1_310 ( .gnd(gnd), .vdd(vdd), .A(_18489_), .B(_17461__bF_buf0), .C(_18490_), .D(_17462__bF_buf0), .Y(_18491_) );
	INVX1 INVX1_2536 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_19_), .Y(_18492_) );
	INVX1 INVX1_2537 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_19_), .Y(_18493_) );
	OAI22X1 OAI22X1_311 ( .gnd(gnd), .vdd(vdd), .A(_18493_), .B(_17467__bF_buf0), .C(_18492_), .D(_17466__bF_buf0), .Y(_18494_) );
	NOR2X1 NOR2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_18491_), .B(_18494_), .Y(_18495_) );
	NAND2X1 NAND2X1_3474 ( .gnd(gnd), .vdd(vdd), .A(_18488_), .B(_18495_), .Y(_18496_) );
	NOR2X1 NOR2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_18481_), .B(_18496_), .Y(_18497_) );
	NAND2X1 NAND2X1_3475 ( .gnd(gnd), .vdd(vdd), .A(_18497_), .B(_18474_), .Y(_428__19_) );
	NAND3X1 NAND3X1_3653 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_20_), .B(_17373__bF_buf3), .C(_17371__bF_buf6), .Y(_18498_) );
	NAND3X1 NAND3X1_3654 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_20_), .B(_17376__bF_buf3), .C(_17371__bF_buf5), .Y(_18499_) );
	NAND2X1 NAND2X1_3476 ( .gnd(gnd), .vdd(vdd), .A(_18498_), .B(_18499_), .Y(_18500_) );
	INVX1 INVX1_2538 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_20_), .Y(_18501_) );
	INVX1 INVX1_2539 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_20_), .Y(_18502_) );
	OAI22X1 OAI22X1_312 ( .gnd(gnd), .vdd(vdd), .A(_18501_), .B(_17384__bF_buf4), .C(_18502_), .D(_17383__bF_buf4), .Y(_18503_) );
	NOR2X1 NOR2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_18500_), .B(_18503_), .Y(_18504_) );
	INVX1 INVX1_2540 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_20_), .Y(_18505_) );
	INVX1 INVX1_2541 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_20_), .Y(_18506_) );
	OAI22X1 OAI22X1_313 ( .gnd(gnd), .vdd(vdd), .A(_18505_), .B(_17394__bF_buf4), .C(_18506_), .D(_17393__bF_buf4), .Y(_18507_) );
	INVX1 INVX1_2542 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_20_), .Y(_18508_) );
	INVX1 INVX1_2543 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_20_), .Y(_18509_) );
	OAI22X1 OAI22X1_314 ( .gnd(gnd), .vdd(vdd), .A(_18508_), .B(_17401__bF_buf4), .C(_18509_), .D(_17400__bF_buf4), .Y(_18510_) );
	NOR2X1 NOR2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_18510_), .B(_18507_), .Y(_18511_) );
	NAND2X1 NAND2X1_3477 ( .gnd(gnd), .vdd(vdd), .A(_18504_), .B(_18511_), .Y(_18512_) );
	INVX1 INVX1_2544 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_20_), .Y(_18513_) );
	INVX1 INVX1_2545 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_20_), .Y(_18514_) );
	OAI22X1 OAI22X1_315 ( .gnd(gnd), .vdd(vdd), .A(_18514_), .B(_17408__bF_buf4), .C(_18513_), .D(_17407__bF_buf4), .Y(_18515_) );
	INVX1 INVX1_2546 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_20_), .Y(_18516_) );
	NAND3X1 NAND3X1_3655 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_20_), .B(_17411__bF_buf5), .C(_17413__bF_buf7), .Y(_18517_) );
	OAI21X1 OAI21X1_3622 ( .gnd(gnd), .vdd(vdd), .A(_18516_), .B(_17412__bF_buf4), .C(_18517_), .Y(_18518_) );
	NOR2X1 NOR2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_18515_), .B(_18518_), .Y(_18519_) );
	INVX1 INVX1_2547 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_20_), .Y(_18520_) );
	NAND3X1 NAND3X1_3656 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(registers_r31_20_), .C(_17419__bF_buf4), .Y(_18521_) );
	OAI21X1 OAI21X1_3623 ( .gnd(gnd), .vdd(vdd), .A(_18520_), .B(_17418__bF_buf4), .C(_18521_), .Y(_18522_) );
	INVX1 INVX1_2548 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_20_), .Y(_18523_) );
	NAND3X1 NAND3X1_3657 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_20_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_18524_) );
	OAI21X1 OAI21X1_3624 ( .gnd(gnd), .vdd(vdd), .A(_18523_), .B(_17423__bF_buf4), .C(_18524_), .Y(_18525_) );
	NOR2X1 NOR2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_18522_), .B(_18525_), .Y(_18526_) );
	NAND2X1 NAND2X1_3478 ( .gnd(gnd), .vdd(vdd), .A(_18526_), .B(_18519_), .Y(_18527_) );
	NOR2X1 NOR2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_18527_), .B(_18512_), .Y(_18528_) );
	AOI22X1 AOI22X1_418 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_20_), .C(registers_r1_20_), .D(_17431__bF_buf4), .Y(_18529_) );
	AOI22X1 AOI22X1_419 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_20_), .C(registers_r5_20_), .D(_17436__bF_buf4), .Y(_18530_) );
	INVX1 INVX1_2549 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_20_), .Y(_18531_) );
	NAND3X1 NAND3X1_3658 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_20_), .B(_17432__bF_buf2), .C(_17392__bF_buf1), .Y(_18532_) );
	OAI21X1 OAI21X1_3625 ( .gnd(gnd), .vdd(vdd), .A(_18531_), .B(_17443__bF_buf4), .C(_18532_), .Y(_18533_) );
	AOI21X1 AOI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_20_), .B(_17440__bF_buf4), .C(_18533_), .Y(_18534_) );
	NAND3X1 NAND3X1_3659 ( .gnd(gnd), .vdd(vdd), .A(_18529_), .B(_18530_), .C(_18534_), .Y(_18535_) );
	INVX1 INVX1_2550 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_20_), .Y(_18536_) );
	INVX1 INVX1_2551 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_20_), .Y(_18537_) );
	OAI22X1 OAI22X1_316 ( .gnd(gnd), .vdd(vdd), .A(_18537_), .B(_17450__bF_buf4), .C(_18536_), .D(_17449__bF_buf4), .Y(_18538_) );
	INVX1 INVX1_2552 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_20_), .Y(_18539_) );
	INVX1 INVX1_2553 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_20_), .Y(_18540_) );
	OAI22X1 OAI22X1_317 ( .gnd(gnd), .vdd(vdd), .A(_18539_), .B(_17456__bF_buf4), .C(_18540_), .D(_17454__bF_buf4), .Y(_18541_) );
	NOR2X1 NOR2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_18541_), .B(_18538_), .Y(_18542_) );
	INVX1 INVX1_2554 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_20_), .Y(_18543_) );
	INVX1 INVX1_2555 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_20_), .Y(_18544_) );
	OAI22X1 OAI22X1_318 ( .gnd(gnd), .vdd(vdd), .A(_18543_), .B(_17461__bF_buf4), .C(_18544_), .D(_17462__bF_buf4), .Y(_18545_) );
	INVX1 INVX1_2556 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_20_), .Y(_18546_) );
	INVX1 INVX1_2557 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_20_), .Y(_18547_) );
	OAI22X1 OAI22X1_319 ( .gnd(gnd), .vdd(vdd), .A(_18547_), .B(_17467__bF_buf4), .C(_18546_), .D(_17466__bF_buf4), .Y(_18548_) );
	NOR2X1 NOR2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_18545_), .B(_18548_), .Y(_18549_) );
	NAND2X1 NAND2X1_3479 ( .gnd(gnd), .vdd(vdd), .A(_18542_), .B(_18549_), .Y(_18550_) );
	NOR2X1 NOR2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_18535_), .B(_18550_), .Y(_18551_) );
	NAND2X1 NAND2X1_3480 ( .gnd(gnd), .vdd(vdd), .A(_18551_), .B(_18528_), .Y(_428__20_) );
	NAND3X1 NAND3X1_3660 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_21_), .B(_17373__bF_buf2), .C(_17371__bF_buf4), .Y(_18552_) );
	NAND3X1 NAND3X1_3661 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_21_), .B(_17376__bF_buf2), .C(_17371__bF_buf3), .Y(_18553_) );
	NAND2X1 NAND2X1_3481 ( .gnd(gnd), .vdd(vdd), .A(_18552_), .B(_18553_), .Y(_18554_) );
	INVX1 INVX1_2558 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_21_), .Y(_18555_) );
	INVX1 INVX1_2559 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_21_), .Y(_18556_) );
	OAI22X1 OAI22X1_320 ( .gnd(gnd), .vdd(vdd), .A(_18555_), .B(_17384__bF_buf3), .C(_18556_), .D(_17383__bF_buf3), .Y(_18557_) );
	NOR2X1 NOR2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_18554_), .B(_18557_), .Y(_18558_) );
	INVX1 INVX1_2560 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_21_), .Y(_18559_) );
	INVX1 INVX1_2561 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_21_), .Y(_18560_) );
	OAI22X1 OAI22X1_321 ( .gnd(gnd), .vdd(vdd), .A(_18559_), .B(_17394__bF_buf3), .C(_18560_), .D(_17393__bF_buf3), .Y(_18561_) );
	INVX1 INVX1_2562 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_21_), .Y(_18562_) );
	INVX1 INVX1_2563 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_21_), .Y(_18563_) );
	OAI22X1 OAI22X1_322 ( .gnd(gnd), .vdd(vdd), .A(_18562_), .B(_17401__bF_buf3), .C(_18563_), .D(_17400__bF_buf3), .Y(_18564_) );
	NOR2X1 NOR2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_18564_), .B(_18561_), .Y(_18565_) );
	NAND2X1 NAND2X1_3482 ( .gnd(gnd), .vdd(vdd), .A(_18558_), .B(_18565_), .Y(_18566_) );
	INVX1 INVX1_2564 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_21_), .Y(_18567_) );
	INVX1 INVX1_2565 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_21_), .Y(_18568_) );
	OAI22X1 OAI22X1_323 ( .gnd(gnd), .vdd(vdd), .A(_18568_), .B(_17408__bF_buf3), .C(_18567_), .D(_17407__bF_buf3), .Y(_18569_) );
	INVX1 INVX1_2566 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_21_), .Y(_18570_) );
	NAND3X1 NAND3X1_3662 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_21_), .B(_17411__bF_buf4), .C(_17413__bF_buf5), .Y(_18571_) );
	OAI21X1 OAI21X1_3626 ( .gnd(gnd), .vdd(vdd), .A(_18570_), .B(_17412__bF_buf3), .C(_18571_), .Y(_18572_) );
	NOR2X1 NOR2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_18569_), .B(_18572_), .Y(_18573_) );
	INVX1 INVX1_2567 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_21_), .Y(_18574_) );
	NAND3X1 NAND3X1_3663 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(registers_r31_21_), .C(_17419__bF_buf3), .Y(_18575_) );
	OAI21X1 OAI21X1_3627 ( .gnd(gnd), .vdd(vdd), .A(_18574_), .B(_17418__bF_buf3), .C(_18575_), .Y(_18576_) );
	INVX1 INVX1_2568 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_21_), .Y(_18577_) );
	NAND3X1 NAND3X1_3664 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_21_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_18578_) );
	OAI21X1 OAI21X1_3628 ( .gnd(gnd), .vdd(vdd), .A(_18577_), .B(_17423__bF_buf3), .C(_18578_), .Y(_18579_) );
	NOR2X1 NOR2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_18576_), .B(_18579_), .Y(_18580_) );
	NAND2X1 NAND2X1_3483 ( .gnd(gnd), .vdd(vdd), .A(_18580_), .B(_18573_), .Y(_18581_) );
	NOR2X1 NOR2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_18581_), .B(_18566_), .Y(_18582_) );
	AOI22X1 AOI22X1_420 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_21_), .C(registers_r1_21_), .D(_17431__bF_buf3), .Y(_18583_) );
	AOI22X1 AOI22X1_421 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_21_), .C(registers_r5_21_), .D(_17436__bF_buf3), .Y(_18584_) );
	INVX1 INVX1_2569 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_21_), .Y(_18585_) );
	NAND3X1 NAND3X1_3665 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_21_), .B(_17432__bF_buf1), .C(_17392__bF_buf7), .Y(_18586_) );
	OAI21X1 OAI21X1_3629 ( .gnd(gnd), .vdd(vdd), .A(_18585_), .B(_17443__bF_buf3), .C(_18586_), .Y(_18587_) );
	AOI21X1 AOI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_21_), .B(_17440__bF_buf3), .C(_18587_), .Y(_18588_) );
	NAND3X1 NAND3X1_3666 ( .gnd(gnd), .vdd(vdd), .A(_18583_), .B(_18584_), .C(_18588_), .Y(_18589_) );
	INVX1 INVX1_2570 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_21_), .Y(_18590_) );
	INVX1 INVX1_2571 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_21_), .Y(_18591_) );
	OAI22X1 OAI22X1_324 ( .gnd(gnd), .vdd(vdd), .A(_18591_), .B(_17450__bF_buf3), .C(_18590_), .D(_17449__bF_buf3), .Y(_18592_) );
	INVX1 INVX1_2572 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_21_), .Y(_18593_) );
	INVX1 INVX1_2573 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_21_), .Y(_18594_) );
	OAI22X1 OAI22X1_325 ( .gnd(gnd), .vdd(vdd), .A(_18593_), .B(_17456__bF_buf3), .C(_18594_), .D(_17454__bF_buf3), .Y(_18595_) );
	NOR2X1 NOR2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_18595_), .B(_18592_), .Y(_18596_) );
	INVX1 INVX1_2574 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_21_), .Y(_18597_) );
	INVX1 INVX1_2575 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_21_), .Y(_18598_) );
	OAI22X1 OAI22X1_326 ( .gnd(gnd), .vdd(vdd), .A(_18597_), .B(_17461__bF_buf3), .C(_18598_), .D(_17462__bF_buf3), .Y(_18599_) );
	INVX1 INVX1_2576 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_21_), .Y(_18600_) );
	INVX1 INVX1_2577 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_21_), .Y(_18601_) );
	OAI22X1 OAI22X1_327 ( .gnd(gnd), .vdd(vdd), .A(_18601_), .B(_17467__bF_buf3), .C(_18600_), .D(_17466__bF_buf3), .Y(_18602_) );
	NOR2X1 NOR2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_18599_), .B(_18602_), .Y(_18603_) );
	NAND2X1 NAND2X1_3484 ( .gnd(gnd), .vdd(vdd), .A(_18596_), .B(_18603_), .Y(_18604_) );
	NOR2X1 NOR2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_18589_), .B(_18604_), .Y(_18605_) );
	NAND2X1 NAND2X1_3485 ( .gnd(gnd), .vdd(vdd), .A(_18605_), .B(_18582_), .Y(_428__21_) );
	NAND3X1 NAND3X1_3667 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_22_), .B(_17373__bF_buf1), .C(_17371__bF_buf2), .Y(_18606_) );
	NAND3X1 NAND3X1_3668 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_22_), .B(_17376__bF_buf1), .C(_17371__bF_buf1), .Y(_18607_) );
	NAND2X1 NAND2X1_3486 ( .gnd(gnd), .vdd(vdd), .A(_18606_), .B(_18607_), .Y(_18608_) );
	INVX1 INVX1_2578 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_22_), .Y(_18609_) );
	INVX1 INVX1_2579 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_22_), .Y(_18610_) );
	OAI22X1 OAI22X1_328 ( .gnd(gnd), .vdd(vdd), .A(_18609_), .B(_17384__bF_buf2), .C(_18610_), .D(_17383__bF_buf2), .Y(_18611_) );
	NOR2X1 NOR2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_18608_), .B(_18611_), .Y(_18612_) );
	INVX1 INVX1_2580 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_22_), .Y(_18613_) );
	INVX1 INVX1_2581 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_22_), .Y(_18614_) );
	OAI22X1 OAI22X1_329 ( .gnd(gnd), .vdd(vdd), .A(_18613_), .B(_17394__bF_buf2), .C(_18614_), .D(_17393__bF_buf2), .Y(_18615_) );
	INVX1 INVX1_2582 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_22_), .Y(_18616_) );
	INVX1 INVX1_2583 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_22_), .Y(_18617_) );
	OAI22X1 OAI22X1_330 ( .gnd(gnd), .vdd(vdd), .A(_18616_), .B(_17401__bF_buf2), .C(_18617_), .D(_17400__bF_buf2), .Y(_18618_) );
	NOR2X1 NOR2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_18618_), .B(_18615_), .Y(_18619_) );
	NAND2X1 NAND2X1_3487 ( .gnd(gnd), .vdd(vdd), .A(_18612_), .B(_18619_), .Y(_18620_) );
	INVX1 INVX1_2584 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_22_), .Y(_18621_) );
	INVX1 INVX1_2585 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_22_), .Y(_18622_) );
	OAI22X1 OAI22X1_331 ( .gnd(gnd), .vdd(vdd), .A(_18622_), .B(_17408__bF_buf2), .C(_18621_), .D(_17407__bF_buf2), .Y(_18623_) );
	INVX1 INVX1_2586 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_22_), .Y(_18624_) );
	NAND3X1 NAND3X1_3669 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_22_), .B(_17411__bF_buf3), .C(_17413__bF_buf3), .Y(_18625_) );
	OAI21X1 OAI21X1_3630 ( .gnd(gnd), .vdd(vdd), .A(_18624_), .B(_17412__bF_buf2), .C(_18625_), .Y(_18626_) );
	NOR2X1 NOR2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_18623_), .B(_18626_), .Y(_18627_) );
	INVX1 INVX1_2587 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_22_), .Y(_18628_) );
	NAND3X1 NAND3X1_3670 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(registers_r31_22_), .C(_17419__bF_buf2), .Y(_18629_) );
	OAI21X1 OAI21X1_3631 ( .gnd(gnd), .vdd(vdd), .A(_18628_), .B(_17418__bF_buf2), .C(_18629_), .Y(_18630_) );
	INVX1 INVX1_2588 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_22_), .Y(_18631_) );
	NAND3X1 NAND3X1_3671 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_22_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_18632_) );
	OAI21X1 OAI21X1_3632 ( .gnd(gnd), .vdd(vdd), .A(_18631_), .B(_17423__bF_buf2), .C(_18632_), .Y(_18633_) );
	NOR2X1 NOR2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_18630_), .B(_18633_), .Y(_18634_) );
	NAND2X1 NAND2X1_3488 ( .gnd(gnd), .vdd(vdd), .A(_18634_), .B(_18627_), .Y(_18635_) );
	NOR2X1 NOR2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_18635_), .B(_18620_), .Y(_18636_) );
	AOI22X1 AOI22X1_422 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf2), .B(registers_a2_22_), .C(registers_r1_22_), .D(_17431__bF_buf2), .Y(_18637_) );
	AOI22X1 AOI22X1_423 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf2), .B(registers_r4_22_), .C(registers_r5_22_), .D(_17436__bF_buf2), .Y(_18638_) );
	INVX1 INVX1_2589 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_22_), .Y(_18639_) );
	NAND3X1 NAND3X1_3672 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_22_), .B(_17432__bF_buf0), .C(_17392__bF_buf5), .Y(_18640_) );
	OAI21X1 OAI21X1_3633 ( .gnd(gnd), .vdd(vdd), .A(_18639_), .B(_17443__bF_buf2), .C(_18640_), .Y(_18641_) );
	AOI21X1 AOI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_22_), .B(_17440__bF_buf2), .C(_18641_), .Y(_18642_) );
	NAND3X1 NAND3X1_3673 ( .gnd(gnd), .vdd(vdd), .A(_18637_), .B(_18638_), .C(_18642_), .Y(_18643_) );
	INVX1 INVX1_2590 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_22_), .Y(_18644_) );
	INVX1 INVX1_2591 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_22_), .Y(_18645_) );
	OAI22X1 OAI22X1_332 ( .gnd(gnd), .vdd(vdd), .A(_18645_), .B(_17450__bF_buf2), .C(_18644_), .D(_17449__bF_buf2), .Y(_18646_) );
	INVX1 INVX1_2592 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_22_), .Y(_18647_) );
	INVX1 INVX1_2593 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_22_), .Y(_18648_) );
	OAI22X1 OAI22X1_333 ( .gnd(gnd), .vdd(vdd), .A(_18647_), .B(_17456__bF_buf2), .C(_18648_), .D(_17454__bF_buf2), .Y(_18649_) );
	NOR2X1 NOR2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_18649_), .B(_18646_), .Y(_18650_) );
	INVX1 INVX1_2594 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_22_), .Y(_18651_) );
	INVX1 INVX1_2595 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_22_), .Y(_18652_) );
	OAI22X1 OAI22X1_334 ( .gnd(gnd), .vdd(vdd), .A(_18651_), .B(_17461__bF_buf2), .C(_18652_), .D(_17462__bF_buf2), .Y(_18653_) );
	INVX1 INVX1_2596 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_22_), .Y(_18654_) );
	INVX1 INVX1_2597 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_22_), .Y(_18655_) );
	OAI22X1 OAI22X1_335 ( .gnd(gnd), .vdd(vdd), .A(_18655_), .B(_17467__bF_buf2), .C(_18654_), .D(_17466__bF_buf2), .Y(_18656_) );
	NOR2X1 NOR2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_18653_), .B(_18656_), .Y(_18657_) );
	NAND2X1 NAND2X1_3489 ( .gnd(gnd), .vdd(vdd), .A(_18650_), .B(_18657_), .Y(_18658_) );
	NOR2X1 NOR2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_18643_), .B(_18658_), .Y(_18659_) );
	NAND2X1 NAND2X1_3490 ( .gnd(gnd), .vdd(vdd), .A(_18659_), .B(_18636_), .Y(_428__22_) );
	NAND3X1 NAND3X1_3674 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_23_), .B(_17373__bF_buf0), .C(_17371__bF_buf0), .Y(_18660_) );
	NAND3X1 NAND3X1_3675 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_23_), .B(_17376__bF_buf0), .C(_17371__bF_buf7), .Y(_18661_) );
	NAND2X1 NAND2X1_3491 ( .gnd(gnd), .vdd(vdd), .A(_18660_), .B(_18661_), .Y(_18662_) );
	INVX1 INVX1_2598 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_23_), .Y(_18663_) );
	INVX1 INVX1_2599 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_23_), .Y(_18664_) );
	OAI22X1 OAI22X1_336 ( .gnd(gnd), .vdd(vdd), .A(_18663_), .B(_17384__bF_buf1), .C(_18664_), .D(_17383__bF_buf1), .Y(_18665_) );
	NOR2X1 NOR2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_18662_), .B(_18665_), .Y(_18666_) );
	INVX1 INVX1_2600 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_23_), .Y(_18667_) );
	INVX1 INVX1_2601 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_23_), .Y(_18668_) );
	OAI22X1 OAI22X1_337 ( .gnd(gnd), .vdd(vdd), .A(_18667_), .B(_17394__bF_buf1), .C(_18668_), .D(_17393__bF_buf1), .Y(_18669_) );
	INVX1 INVX1_2602 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_23_), .Y(_18670_) );
	INVX1 INVX1_2603 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_23_), .Y(_18671_) );
	OAI22X1 OAI22X1_338 ( .gnd(gnd), .vdd(vdd), .A(_18670_), .B(_17401__bF_buf1), .C(_18671_), .D(_17400__bF_buf1), .Y(_18672_) );
	NOR2X1 NOR2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_18672_), .B(_18669_), .Y(_18673_) );
	NAND2X1 NAND2X1_3492 ( .gnd(gnd), .vdd(vdd), .A(_18666_), .B(_18673_), .Y(_18674_) );
	INVX1 INVX1_2604 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_23_), .Y(_18675_) );
	INVX1 INVX1_2605 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_23_), .Y(_18676_) );
	OAI22X1 OAI22X1_339 ( .gnd(gnd), .vdd(vdd), .A(_18676_), .B(_17408__bF_buf1), .C(_18675_), .D(_17407__bF_buf1), .Y(_18677_) );
	INVX1 INVX1_2606 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_23_), .Y(_18678_) );
	NAND3X1 NAND3X1_3676 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_23_), .B(_17411__bF_buf2), .C(_17413__bF_buf1), .Y(_18679_) );
	OAI21X1 OAI21X1_3634 ( .gnd(gnd), .vdd(vdd), .A(_18678_), .B(_17412__bF_buf1), .C(_18679_), .Y(_18680_) );
	NOR2X1 NOR2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_18677_), .B(_18680_), .Y(_18681_) );
	INVX1 INVX1_2607 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_23_), .Y(_18682_) );
	NAND3X1 NAND3X1_3677 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(registers_r31_23_), .C(_17419__bF_buf1), .Y(_18683_) );
	OAI21X1 OAI21X1_3635 ( .gnd(gnd), .vdd(vdd), .A(_18682_), .B(_17418__bF_buf1), .C(_18683_), .Y(_18684_) );
	INVX1 INVX1_2608 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_23_), .Y(_18685_) );
	NAND3X1 NAND3X1_3678 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_23_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_18686_) );
	OAI21X1 OAI21X1_3636 ( .gnd(gnd), .vdd(vdd), .A(_18685_), .B(_17423__bF_buf1), .C(_18686_), .Y(_18687_) );
	NOR2X1 NOR2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_18684_), .B(_18687_), .Y(_18688_) );
	NAND2X1 NAND2X1_3493 ( .gnd(gnd), .vdd(vdd), .A(_18688_), .B(_18681_), .Y(_18689_) );
	NOR2X1 NOR2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_18689_), .B(_18674_), .Y(_18690_) );
	AOI22X1 AOI22X1_424 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf1), .B(registers_a2_23_), .C(registers_r1_23_), .D(_17431__bF_buf1), .Y(_18691_) );
	AOI22X1 AOI22X1_425 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf1), .B(registers_r4_23_), .C(registers_r5_23_), .D(_17436__bF_buf1), .Y(_18692_) );
	INVX1 INVX1_2609 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_23_), .Y(_18693_) );
	NAND3X1 NAND3X1_3679 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_23_), .B(_17432__bF_buf4), .C(_17392__bF_buf3), .Y(_18694_) );
	OAI21X1 OAI21X1_3637 ( .gnd(gnd), .vdd(vdd), .A(_18693_), .B(_17443__bF_buf1), .C(_18694_), .Y(_18695_) );
	AOI21X1 AOI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_23_), .B(_17440__bF_buf1), .C(_18695_), .Y(_18696_) );
	NAND3X1 NAND3X1_3680 ( .gnd(gnd), .vdd(vdd), .A(_18691_), .B(_18692_), .C(_18696_), .Y(_18697_) );
	INVX1 INVX1_2610 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_23_), .Y(_18698_) );
	INVX1 INVX1_2611 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_23_), .Y(_18699_) );
	OAI22X1 OAI22X1_340 ( .gnd(gnd), .vdd(vdd), .A(_18699_), .B(_17450__bF_buf1), .C(_18698_), .D(_17449__bF_buf1), .Y(_18700_) );
	INVX1 INVX1_2612 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_23_), .Y(_18701_) );
	INVX1 INVX1_2613 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_23_), .Y(_18702_) );
	OAI22X1 OAI22X1_341 ( .gnd(gnd), .vdd(vdd), .A(_18701_), .B(_17456__bF_buf1), .C(_18702_), .D(_17454__bF_buf1), .Y(_18703_) );
	NOR2X1 NOR2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_18703_), .B(_18700_), .Y(_18704_) );
	INVX1 INVX1_2614 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_23_), .Y(_18705_) );
	INVX1 INVX1_2615 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_23_), .Y(_18706_) );
	OAI22X1 OAI22X1_342 ( .gnd(gnd), .vdd(vdd), .A(_18705_), .B(_17461__bF_buf1), .C(_18706_), .D(_17462__bF_buf1), .Y(_18707_) );
	INVX1 INVX1_2616 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_23_), .Y(_18708_) );
	INVX1 INVX1_2617 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_23_), .Y(_18709_) );
	OAI22X1 OAI22X1_343 ( .gnd(gnd), .vdd(vdd), .A(_18709_), .B(_17467__bF_buf1), .C(_18708_), .D(_17466__bF_buf1), .Y(_18710_) );
	NOR2X1 NOR2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_18707_), .B(_18710_), .Y(_18711_) );
	NAND2X1 NAND2X1_3494 ( .gnd(gnd), .vdd(vdd), .A(_18704_), .B(_18711_), .Y(_18712_) );
	NOR2X1 NOR2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_18697_), .B(_18712_), .Y(_18713_) );
	NAND2X1 NAND2X1_3495 ( .gnd(gnd), .vdd(vdd), .A(_18713_), .B(_18690_), .Y(_428__23_) );
	NAND3X1 NAND3X1_3681 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_24_), .B(_17373__bF_buf5), .C(_17371__bF_buf6), .Y(_18714_) );
	NAND3X1 NAND3X1_3682 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_24_), .B(_17376__bF_buf5), .C(_17371__bF_buf5), .Y(_18715_) );
	NAND2X1 NAND2X1_3496 ( .gnd(gnd), .vdd(vdd), .A(_18714_), .B(_18715_), .Y(_18716_) );
	INVX1 INVX1_2618 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_24_), .Y(_18717_) );
	INVX1 INVX1_2619 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_24_), .Y(_18718_) );
	OAI22X1 OAI22X1_344 ( .gnd(gnd), .vdd(vdd), .A(_18717_), .B(_17384__bF_buf0), .C(_18718_), .D(_17383__bF_buf0), .Y(_18719_) );
	NOR2X1 NOR2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_18716_), .B(_18719_), .Y(_18720_) );
	INVX1 INVX1_2620 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_24_), .Y(_18721_) );
	INVX1 INVX1_2621 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_24_), .Y(_18722_) );
	OAI22X1 OAI22X1_345 ( .gnd(gnd), .vdd(vdd), .A(_18721_), .B(_17394__bF_buf0), .C(_18722_), .D(_17393__bF_buf0), .Y(_18723_) );
	INVX1 INVX1_2622 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_24_), .Y(_18724_) );
	INVX1 INVX1_2623 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_24_), .Y(_18725_) );
	OAI22X1 OAI22X1_346 ( .gnd(gnd), .vdd(vdd), .A(_18724_), .B(_17401__bF_buf0), .C(_18725_), .D(_17400__bF_buf0), .Y(_18726_) );
	NOR2X1 NOR2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_18726_), .B(_18723_), .Y(_18727_) );
	NAND2X1 NAND2X1_3497 ( .gnd(gnd), .vdd(vdd), .A(_18720_), .B(_18727_), .Y(_18728_) );
	INVX1 INVX1_2624 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_24_), .Y(_18729_) );
	INVX1 INVX1_2625 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_24_), .Y(_18730_) );
	OAI22X1 OAI22X1_347 ( .gnd(gnd), .vdd(vdd), .A(_18730_), .B(_17408__bF_buf0), .C(_18729_), .D(_17407__bF_buf0), .Y(_18731_) );
	INVX1 INVX1_2626 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_24_), .Y(_18732_) );
	NAND3X1 NAND3X1_3683 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_24_), .B(_17411__bF_buf1), .C(_17413__bF_buf7), .Y(_18733_) );
	OAI21X1 OAI21X1_3638 ( .gnd(gnd), .vdd(vdd), .A(_18732_), .B(_17412__bF_buf0), .C(_18733_), .Y(_18734_) );
	NOR2X1 NOR2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_18731_), .B(_18734_), .Y(_18735_) );
	INVX1 INVX1_2627 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_24_), .Y(_18736_) );
	NAND3X1 NAND3X1_3684 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(registers_r31_24_), .C(_17419__bF_buf0), .Y(_18737_) );
	OAI21X1 OAI21X1_3639 ( .gnd(gnd), .vdd(vdd), .A(_18736_), .B(_17418__bF_buf0), .C(_18737_), .Y(_18738_) );
	INVX1 INVX1_2628 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_24_), .Y(_18739_) );
	NAND3X1 NAND3X1_3685 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_24_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_18740_) );
	OAI21X1 OAI21X1_3640 ( .gnd(gnd), .vdd(vdd), .A(_18739_), .B(_17423__bF_buf0), .C(_18740_), .Y(_18741_) );
	NOR2X1 NOR2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_18738_), .B(_18741_), .Y(_18742_) );
	NAND2X1 NAND2X1_3498 ( .gnd(gnd), .vdd(vdd), .A(_18742_), .B(_18735_), .Y(_18743_) );
	NOR2X1 NOR2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_18743_), .B(_18728_), .Y(_18744_) );
	AOI22X1 AOI22X1_426 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf0), .B(registers_a2_24_), .C(registers_r1_24_), .D(_17431__bF_buf0), .Y(_18745_) );
	AOI22X1 AOI22X1_427 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf0), .B(registers_r4_24_), .C(registers_r5_24_), .D(_17436__bF_buf0), .Y(_18746_) );
	INVX1 INVX1_2629 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_24_), .Y(_18747_) );
	NAND3X1 NAND3X1_3686 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_24_), .B(_17432__bF_buf3), .C(_17392__bF_buf1), .Y(_18748_) );
	OAI21X1 OAI21X1_3641 ( .gnd(gnd), .vdd(vdd), .A(_18747_), .B(_17443__bF_buf0), .C(_18748_), .Y(_18749_) );
	AOI21X1 AOI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_24_), .B(_17440__bF_buf0), .C(_18749_), .Y(_18750_) );
	NAND3X1 NAND3X1_3687 ( .gnd(gnd), .vdd(vdd), .A(_18745_), .B(_18746_), .C(_18750_), .Y(_18751_) );
	INVX1 INVX1_2630 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_24_), .Y(_18752_) );
	INVX1 INVX1_2631 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_24_), .Y(_18753_) );
	OAI22X1 OAI22X1_348 ( .gnd(gnd), .vdd(vdd), .A(_18753_), .B(_17450__bF_buf0), .C(_18752_), .D(_17449__bF_buf0), .Y(_18754_) );
	INVX1 INVX1_2632 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_24_), .Y(_18755_) );
	INVX1 INVX1_2633 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_24_), .Y(_18756_) );
	OAI22X1 OAI22X1_349 ( .gnd(gnd), .vdd(vdd), .A(_18755_), .B(_17456__bF_buf0), .C(_18756_), .D(_17454__bF_buf0), .Y(_18757_) );
	NOR2X1 NOR2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_18757_), .B(_18754_), .Y(_18758_) );
	INVX1 INVX1_2634 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_24_), .Y(_18759_) );
	INVX1 INVX1_2635 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_24_), .Y(_18760_) );
	OAI22X1 OAI22X1_350 ( .gnd(gnd), .vdd(vdd), .A(_18759_), .B(_17461__bF_buf0), .C(_18760_), .D(_17462__bF_buf0), .Y(_18761_) );
	INVX1 INVX1_2636 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_24_), .Y(_18762_) );
	INVX1 INVX1_2637 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_24_), .Y(_18763_) );
	OAI22X1 OAI22X1_351 ( .gnd(gnd), .vdd(vdd), .A(_18763_), .B(_17467__bF_buf0), .C(_18762_), .D(_17466__bF_buf0), .Y(_18764_) );
	NOR2X1 NOR2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_18761_), .B(_18764_), .Y(_18765_) );
	NAND2X1 NAND2X1_3499 ( .gnd(gnd), .vdd(vdd), .A(_18758_), .B(_18765_), .Y(_18766_) );
	NOR2X1 NOR2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_18751_), .B(_18766_), .Y(_18767_) );
	NAND2X1 NAND2X1_3500 ( .gnd(gnd), .vdd(vdd), .A(_18767_), .B(_18744_), .Y(_428__24_) );
	NAND3X1 NAND3X1_3688 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_25_), .B(_17373__bF_buf4), .C(_17371__bF_buf4), .Y(_18768_) );
	NAND3X1 NAND3X1_3689 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_25_), .B(_17376__bF_buf4), .C(_17371__bF_buf3), .Y(_18769_) );
	NAND2X1 NAND2X1_3501 ( .gnd(gnd), .vdd(vdd), .A(_18768_), .B(_18769_), .Y(_18770_) );
	INVX1 INVX1_2638 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_25_), .Y(_18771_) );
	INVX1 INVX1_2639 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_25_), .Y(_18772_) );
	OAI22X1 OAI22X1_352 ( .gnd(gnd), .vdd(vdd), .A(_18771_), .B(_17384__bF_buf4), .C(_18772_), .D(_17383__bF_buf4), .Y(_18773_) );
	NOR2X1 NOR2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_18770_), .B(_18773_), .Y(_18774_) );
	INVX1 INVX1_2640 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_25_), .Y(_18775_) );
	INVX1 INVX1_2641 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_25_), .Y(_18776_) );
	OAI22X1 OAI22X1_353 ( .gnd(gnd), .vdd(vdd), .A(_18775_), .B(_17394__bF_buf4), .C(_18776_), .D(_17393__bF_buf4), .Y(_18777_) );
	INVX1 INVX1_2642 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_25_), .Y(_18778_) );
	INVX1 INVX1_2643 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_25_), .Y(_18779_) );
	OAI22X1 OAI22X1_354 ( .gnd(gnd), .vdd(vdd), .A(_18778_), .B(_17401__bF_buf4), .C(_18779_), .D(_17400__bF_buf4), .Y(_18780_) );
	NOR2X1 NOR2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_18780_), .B(_18777_), .Y(_18781_) );
	NAND2X1 NAND2X1_3502 ( .gnd(gnd), .vdd(vdd), .A(_18774_), .B(_18781_), .Y(_18782_) );
	INVX1 INVX1_2644 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_25_), .Y(_18783_) );
	INVX1 INVX1_2645 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_25_), .Y(_18784_) );
	OAI22X1 OAI22X1_355 ( .gnd(gnd), .vdd(vdd), .A(_18784_), .B(_17408__bF_buf4), .C(_18783_), .D(_17407__bF_buf4), .Y(_18785_) );
	INVX1 INVX1_2646 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_25_), .Y(_18786_) );
	NAND3X1 NAND3X1_3690 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_25_), .B(_17411__bF_buf0), .C(_17413__bF_buf5), .Y(_18787_) );
	OAI21X1 OAI21X1_3642 ( .gnd(gnd), .vdd(vdd), .A(_18786_), .B(_17412__bF_buf4), .C(_18787_), .Y(_18788_) );
	NOR2X1 NOR2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_18785_), .B(_18788_), .Y(_18789_) );
	INVX1 INVX1_2647 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_25_), .Y(_18790_) );
	NAND3X1 NAND3X1_3691 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf4), .B(registers_r31_25_), .C(_17419__bF_buf4), .Y(_18791_) );
	OAI21X1 OAI21X1_3643 ( .gnd(gnd), .vdd(vdd), .A(_18790_), .B(_17418__bF_buf4), .C(_18791_), .Y(_18792_) );
	INVX1 INVX1_2648 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_25_), .Y(_18793_) );
	NAND3X1 NAND3X1_3692 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_25_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_18794_) );
	OAI21X1 OAI21X1_3644 ( .gnd(gnd), .vdd(vdd), .A(_18793_), .B(_17423__bF_buf4), .C(_18794_), .Y(_18795_) );
	NOR2X1 NOR2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_18792_), .B(_18795_), .Y(_18796_) );
	NAND2X1 NAND2X1_3503 ( .gnd(gnd), .vdd(vdd), .A(_18796_), .B(_18789_), .Y(_18797_) );
	NOR2X1 NOR2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_18797_), .B(_18782_), .Y(_18798_) );
	AOI22X1 AOI22X1_428 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_25_), .C(registers_r1_25_), .D(_17431__bF_buf4), .Y(_18799_) );
	AOI22X1 AOI22X1_429 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_25_), .C(registers_r5_25_), .D(_17436__bF_buf4), .Y(_18800_) );
	INVX1 INVX1_2649 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_25_), .Y(_18801_) );
	NAND3X1 NAND3X1_3693 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_25_), .B(_17432__bF_buf2), .C(_17392__bF_buf7), .Y(_18802_) );
	OAI21X1 OAI21X1_3645 ( .gnd(gnd), .vdd(vdd), .A(_18801_), .B(_17443__bF_buf4), .C(_18802_), .Y(_18803_) );
	AOI21X1 AOI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_25_), .B(_17440__bF_buf4), .C(_18803_), .Y(_18804_) );
	NAND3X1 NAND3X1_3694 ( .gnd(gnd), .vdd(vdd), .A(_18799_), .B(_18800_), .C(_18804_), .Y(_18805_) );
	INVX1 INVX1_2650 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_25_), .Y(_18806_) );
	INVX1 INVX1_2651 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_25_), .Y(_18807_) );
	OAI22X1 OAI22X1_356 ( .gnd(gnd), .vdd(vdd), .A(_18807_), .B(_17450__bF_buf4), .C(_18806_), .D(_17449__bF_buf4), .Y(_18808_) );
	INVX1 INVX1_2652 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_25_), .Y(_18809_) );
	INVX1 INVX1_2653 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_25_), .Y(_18810_) );
	OAI22X1 OAI22X1_357 ( .gnd(gnd), .vdd(vdd), .A(_18809_), .B(_17456__bF_buf4), .C(_18810_), .D(_17454__bF_buf4), .Y(_18811_) );
	NOR2X1 NOR2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_18811_), .B(_18808_), .Y(_18812_) );
	INVX1 INVX1_2654 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_25_), .Y(_18813_) );
	INVX1 INVX1_2655 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_25_), .Y(_18814_) );
	OAI22X1 OAI22X1_358 ( .gnd(gnd), .vdd(vdd), .A(_18813_), .B(_17461__bF_buf4), .C(_18814_), .D(_17462__bF_buf4), .Y(_18815_) );
	INVX1 INVX1_2656 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_25_), .Y(_18816_) );
	INVX1 INVX1_2657 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_25_), .Y(_18817_) );
	OAI22X1 OAI22X1_359 ( .gnd(gnd), .vdd(vdd), .A(_18817_), .B(_17467__bF_buf4), .C(_18816_), .D(_17466__bF_buf4), .Y(_18818_) );
	NOR2X1 NOR2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_18815_), .B(_18818_), .Y(_18819_) );
	NAND2X1 NAND2X1_3504 ( .gnd(gnd), .vdd(vdd), .A(_18812_), .B(_18819_), .Y(_18820_) );
	NOR2X1 NOR2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_18805_), .B(_18820_), .Y(_18821_) );
	NAND2X1 NAND2X1_3505 ( .gnd(gnd), .vdd(vdd), .A(_18821_), .B(_18798_), .Y(_428__25_) );
	NAND3X1 NAND3X1_3695 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_26_), .B(_17373__bF_buf3), .C(_17371__bF_buf2), .Y(_18822_) );
	NAND3X1 NAND3X1_3696 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_26_), .B(_17376__bF_buf3), .C(_17371__bF_buf1), .Y(_18823_) );
	NAND2X1 NAND2X1_3506 ( .gnd(gnd), .vdd(vdd), .A(_18822_), .B(_18823_), .Y(_18824_) );
	INVX1 INVX1_2658 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_26_), .Y(_18825_) );
	INVX1 INVX1_2659 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_26_), .Y(_18826_) );
	OAI22X1 OAI22X1_360 ( .gnd(gnd), .vdd(vdd), .A(_18825_), .B(_17384__bF_buf3), .C(_18826_), .D(_17383__bF_buf3), .Y(_18827_) );
	NOR2X1 NOR2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_18824_), .B(_18827_), .Y(_18828_) );
	INVX1 INVX1_2660 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_26_), .Y(_18829_) );
	INVX1 INVX1_2661 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_26_), .Y(_18830_) );
	OAI22X1 OAI22X1_361 ( .gnd(gnd), .vdd(vdd), .A(_18829_), .B(_17394__bF_buf3), .C(_18830_), .D(_17393__bF_buf3), .Y(_18831_) );
	INVX1 INVX1_2662 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_26_), .Y(_18832_) );
	INVX1 INVX1_2663 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_26_), .Y(_18833_) );
	OAI22X1 OAI22X1_362 ( .gnd(gnd), .vdd(vdd), .A(_18832_), .B(_17401__bF_buf3), .C(_18833_), .D(_17400__bF_buf3), .Y(_18834_) );
	NOR2X1 NOR2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_18834_), .B(_18831_), .Y(_18835_) );
	NAND2X1 NAND2X1_3507 ( .gnd(gnd), .vdd(vdd), .A(_18828_), .B(_18835_), .Y(_18836_) );
	INVX1 INVX1_2664 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_26_), .Y(_18837_) );
	INVX1 INVX1_2665 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_26_), .Y(_18838_) );
	OAI22X1 OAI22X1_363 ( .gnd(gnd), .vdd(vdd), .A(_18838_), .B(_17408__bF_buf3), .C(_18837_), .D(_17407__bF_buf3), .Y(_18839_) );
	INVX1 INVX1_2666 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_26_), .Y(_18840_) );
	NAND3X1 NAND3X1_3697 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_26_), .B(_17411__bF_buf5), .C(_17413__bF_buf3), .Y(_18841_) );
	OAI21X1 OAI21X1_3646 ( .gnd(gnd), .vdd(vdd), .A(_18840_), .B(_17412__bF_buf3), .C(_18841_), .Y(_18842_) );
	NOR2X1 NOR2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_18839_), .B(_18842_), .Y(_18843_) );
	INVX1 INVX1_2667 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_26_), .Y(_18844_) );
	NAND3X1 NAND3X1_3698 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf3), .B(registers_r31_26_), .C(_17419__bF_buf3), .Y(_18845_) );
	OAI21X1 OAI21X1_3647 ( .gnd(gnd), .vdd(vdd), .A(_18844_), .B(_17418__bF_buf3), .C(_18845_), .Y(_18846_) );
	INVX1 INVX1_2668 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_26_), .Y(_18847_) );
	NAND3X1 NAND3X1_3699 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_26_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_18848_) );
	OAI21X1 OAI21X1_3648 ( .gnd(gnd), .vdd(vdd), .A(_18847_), .B(_17423__bF_buf3), .C(_18848_), .Y(_18849_) );
	NOR2X1 NOR2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_18846_), .B(_18849_), .Y(_18850_) );
	NAND2X1 NAND2X1_3508 ( .gnd(gnd), .vdd(vdd), .A(_18850_), .B(_18843_), .Y(_18851_) );
	NOR2X1 NOR2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_18851_), .B(_18836_), .Y(_18852_) );
	AOI22X1 AOI22X1_430 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_26_), .C(registers_r1_26_), .D(_17431__bF_buf3), .Y(_18853_) );
	AOI22X1 AOI22X1_431 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_26_), .C(registers_r5_26_), .D(_17436__bF_buf3), .Y(_18854_) );
	INVX1 INVX1_2669 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_26_), .Y(_18855_) );
	NAND3X1 NAND3X1_3700 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_26_), .B(_17432__bF_buf1), .C(_17392__bF_buf5), .Y(_18856_) );
	OAI21X1 OAI21X1_3649 ( .gnd(gnd), .vdd(vdd), .A(_18855_), .B(_17443__bF_buf3), .C(_18856_), .Y(_18857_) );
	AOI21X1 AOI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_26_), .B(_17440__bF_buf3), .C(_18857_), .Y(_18858_) );
	NAND3X1 NAND3X1_3701 ( .gnd(gnd), .vdd(vdd), .A(_18853_), .B(_18854_), .C(_18858_), .Y(_18859_) );
	INVX1 INVX1_2670 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_26_), .Y(_18860_) );
	INVX1 INVX1_2671 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_26_), .Y(_18861_) );
	OAI22X1 OAI22X1_364 ( .gnd(gnd), .vdd(vdd), .A(_18861_), .B(_17450__bF_buf3), .C(_18860_), .D(_17449__bF_buf3), .Y(_18862_) );
	INVX1 INVX1_2672 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_26_), .Y(_18863_) );
	INVX1 INVX1_2673 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_26_), .Y(_18864_) );
	OAI22X1 OAI22X1_365 ( .gnd(gnd), .vdd(vdd), .A(_18863_), .B(_17456__bF_buf3), .C(_18864_), .D(_17454__bF_buf3), .Y(_18865_) );
	NOR2X1 NOR2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_18865_), .B(_18862_), .Y(_18866_) );
	INVX1 INVX1_2674 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_26_), .Y(_18867_) );
	INVX1 INVX1_2675 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_26_), .Y(_18868_) );
	OAI22X1 OAI22X1_366 ( .gnd(gnd), .vdd(vdd), .A(_18867_), .B(_17461__bF_buf3), .C(_18868_), .D(_17462__bF_buf3), .Y(_18869_) );
	INVX1 INVX1_2676 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_26_), .Y(_18870_) );
	INVX1 INVX1_2677 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_26_), .Y(_18871_) );
	OAI22X1 OAI22X1_367 ( .gnd(gnd), .vdd(vdd), .A(_18871_), .B(_17467__bF_buf3), .C(_18870_), .D(_17466__bF_buf3), .Y(_18872_) );
	NOR2X1 NOR2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_18869_), .B(_18872_), .Y(_18873_) );
	NAND2X1 NAND2X1_3509 ( .gnd(gnd), .vdd(vdd), .A(_18866_), .B(_18873_), .Y(_18874_) );
	NOR2X1 NOR2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_18859_), .B(_18874_), .Y(_18875_) );
	NAND2X1 NAND2X1_3510 ( .gnd(gnd), .vdd(vdd), .A(_18875_), .B(_18852_), .Y(_428__26_) );
	NAND3X1 NAND3X1_3702 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_27_), .B(_17373__bF_buf2), .C(_17371__bF_buf0), .Y(_18876_) );
	NAND3X1 NAND3X1_3703 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_27_), .B(_17376__bF_buf2), .C(_17371__bF_buf7), .Y(_18877_) );
	NAND2X1 NAND2X1_3511 ( .gnd(gnd), .vdd(vdd), .A(_18876_), .B(_18877_), .Y(_18878_) );
	INVX1 INVX1_2678 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_27_), .Y(_18879_) );
	INVX1 INVX1_2679 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_27_), .Y(_18880_) );
	OAI22X1 OAI22X1_368 ( .gnd(gnd), .vdd(vdd), .A(_18879_), .B(_17384__bF_buf2), .C(_18880_), .D(_17383__bF_buf2), .Y(_18881_) );
	NOR2X1 NOR2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_18878_), .B(_18881_), .Y(_18882_) );
	INVX1 INVX1_2680 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_27_), .Y(_18883_) );
	INVX1 INVX1_2681 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_27_), .Y(_18884_) );
	OAI22X1 OAI22X1_369 ( .gnd(gnd), .vdd(vdd), .A(_18883_), .B(_17394__bF_buf2), .C(_18884_), .D(_17393__bF_buf2), .Y(_18885_) );
	INVX1 INVX1_2682 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_27_), .Y(_18886_) );
	INVX1 INVX1_2683 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_27_), .Y(_18887_) );
	OAI22X1 OAI22X1_370 ( .gnd(gnd), .vdd(vdd), .A(_18886_), .B(_17401__bF_buf2), .C(_18887_), .D(_17400__bF_buf2), .Y(_18888_) );
	NOR2X1 NOR2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_18888_), .B(_18885_), .Y(_18889_) );
	NAND2X1 NAND2X1_3512 ( .gnd(gnd), .vdd(vdd), .A(_18882_), .B(_18889_), .Y(_18890_) );
	INVX1 INVX1_2684 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_27_), .Y(_18891_) );
	INVX1 INVX1_2685 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_27_), .Y(_18892_) );
	OAI22X1 OAI22X1_371 ( .gnd(gnd), .vdd(vdd), .A(_18892_), .B(_17408__bF_buf2), .C(_18891_), .D(_17407__bF_buf2), .Y(_18893_) );
	INVX1 INVX1_2686 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_27_), .Y(_18894_) );
	NAND3X1 NAND3X1_3704 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_27_), .B(_17411__bF_buf4), .C(_17413__bF_buf1), .Y(_18895_) );
	OAI21X1 OAI21X1_3650 ( .gnd(gnd), .vdd(vdd), .A(_18894_), .B(_17412__bF_buf2), .C(_18895_), .Y(_18896_) );
	NOR2X1 NOR2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_18893_), .B(_18896_), .Y(_18897_) );
	INVX1 INVX1_2687 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_27_), .Y(_18898_) );
	NAND3X1 NAND3X1_3705 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf2), .B(registers_r31_27_), .C(_17419__bF_buf2), .Y(_18899_) );
	OAI21X1 OAI21X1_3651 ( .gnd(gnd), .vdd(vdd), .A(_18898_), .B(_17418__bF_buf2), .C(_18899_), .Y(_18900_) );
	INVX1 INVX1_2688 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_27_), .Y(_18901_) );
	NAND3X1 NAND3X1_3706 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_27_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_18902_) );
	OAI21X1 OAI21X1_3652 ( .gnd(gnd), .vdd(vdd), .A(_18901_), .B(_17423__bF_buf2), .C(_18902_), .Y(_18903_) );
	NOR2X1 NOR2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_18900_), .B(_18903_), .Y(_18904_) );
	NAND2X1 NAND2X1_3513 ( .gnd(gnd), .vdd(vdd), .A(_18904_), .B(_18897_), .Y(_18905_) );
	NOR2X1 NOR2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_18905_), .B(_18890_), .Y(_18906_) );
	AOI22X1 AOI22X1_432 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf2), .B(registers_a2_27_), .C(registers_r1_27_), .D(_17431__bF_buf2), .Y(_18907_) );
	AOI22X1 AOI22X1_433 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf2), .B(registers_r4_27_), .C(registers_r5_27_), .D(_17436__bF_buf2), .Y(_18908_) );
	INVX1 INVX1_2689 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_27_), .Y(_18909_) );
	NAND3X1 NAND3X1_3707 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_27_), .B(_17432__bF_buf0), .C(_17392__bF_buf3), .Y(_18910_) );
	OAI21X1 OAI21X1_3653 ( .gnd(gnd), .vdd(vdd), .A(_18909_), .B(_17443__bF_buf2), .C(_18910_), .Y(_18911_) );
	AOI21X1 AOI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_27_), .B(_17440__bF_buf2), .C(_18911_), .Y(_18912_) );
	NAND3X1 NAND3X1_3708 ( .gnd(gnd), .vdd(vdd), .A(_18907_), .B(_18908_), .C(_18912_), .Y(_18913_) );
	INVX1 INVX1_2690 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_27_), .Y(_18914_) );
	INVX1 INVX1_2691 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_27_), .Y(_18915_) );
	OAI22X1 OAI22X1_372 ( .gnd(gnd), .vdd(vdd), .A(_18915_), .B(_17450__bF_buf2), .C(_18914_), .D(_17449__bF_buf2), .Y(_18916_) );
	INVX1 INVX1_2692 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_27_), .Y(_18917_) );
	INVX1 INVX1_2693 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_27_), .Y(_18918_) );
	OAI22X1 OAI22X1_373 ( .gnd(gnd), .vdd(vdd), .A(_18917_), .B(_17456__bF_buf2), .C(_18918_), .D(_17454__bF_buf2), .Y(_18919_) );
	NOR2X1 NOR2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_18919_), .B(_18916_), .Y(_18920_) );
	INVX1 INVX1_2694 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_27_), .Y(_18921_) );
	INVX1 INVX1_2695 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_27_), .Y(_18922_) );
	OAI22X1 OAI22X1_374 ( .gnd(gnd), .vdd(vdd), .A(_18921_), .B(_17461__bF_buf2), .C(_18922_), .D(_17462__bF_buf2), .Y(_18923_) );
	INVX1 INVX1_2696 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_27_), .Y(_18924_) );
	INVX1 INVX1_2697 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_27_), .Y(_18925_) );
	OAI22X1 OAI22X1_375 ( .gnd(gnd), .vdd(vdd), .A(_18925_), .B(_17467__bF_buf2), .C(_18924_), .D(_17466__bF_buf2), .Y(_18926_) );
	NOR2X1 NOR2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_18923_), .B(_18926_), .Y(_18927_) );
	NAND2X1 NAND2X1_3514 ( .gnd(gnd), .vdd(vdd), .A(_18920_), .B(_18927_), .Y(_18928_) );
	NOR2X1 NOR2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_18913_), .B(_18928_), .Y(_18929_) );
	NAND2X1 NAND2X1_3515 ( .gnd(gnd), .vdd(vdd), .A(_18929_), .B(_18906_), .Y(_428__27_) );
	NAND3X1 NAND3X1_3709 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_28_), .B(_17373__bF_buf1), .C(_17371__bF_buf6), .Y(_18930_) );
	NAND3X1 NAND3X1_3710 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_28_), .B(_17376__bF_buf1), .C(_17371__bF_buf5), .Y(_18931_) );
	NAND2X1 NAND2X1_3516 ( .gnd(gnd), .vdd(vdd), .A(_18930_), .B(_18931_), .Y(_18932_) );
	INVX1 INVX1_2698 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_28_), .Y(_18933_) );
	INVX1 INVX1_2699 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_28_), .Y(_18934_) );
	OAI22X1 OAI22X1_376 ( .gnd(gnd), .vdd(vdd), .A(_18933_), .B(_17384__bF_buf1), .C(_18934_), .D(_17383__bF_buf1), .Y(_18935_) );
	NOR2X1 NOR2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_18932_), .B(_18935_), .Y(_18936_) );
	INVX1 INVX1_2700 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_28_), .Y(_18937_) );
	INVX1 INVX1_2701 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_28_), .Y(_18938_) );
	OAI22X1 OAI22X1_377 ( .gnd(gnd), .vdd(vdd), .A(_18937_), .B(_17394__bF_buf1), .C(_18938_), .D(_17393__bF_buf1), .Y(_18939_) );
	INVX1 INVX1_2702 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_28_), .Y(_18940_) );
	INVX1 INVX1_2703 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_28_), .Y(_18941_) );
	OAI22X1 OAI22X1_378 ( .gnd(gnd), .vdd(vdd), .A(_18940_), .B(_17401__bF_buf1), .C(_18941_), .D(_17400__bF_buf1), .Y(_18942_) );
	NOR2X1 NOR2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_18942_), .B(_18939_), .Y(_18943_) );
	NAND2X1 NAND2X1_3517 ( .gnd(gnd), .vdd(vdd), .A(_18936_), .B(_18943_), .Y(_18944_) );
	INVX1 INVX1_2704 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_28_), .Y(_18945_) );
	INVX1 INVX1_2705 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_28_), .Y(_18946_) );
	OAI22X1 OAI22X1_379 ( .gnd(gnd), .vdd(vdd), .A(_18946_), .B(_17408__bF_buf1), .C(_18945_), .D(_17407__bF_buf1), .Y(_18947_) );
	INVX1 INVX1_2706 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_28_), .Y(_18948_) );
	NAND3X1 NAND3X1_3711 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_28_), .B(_17411__bF_buf3), .C(_17413__bF_buf7), .Y(_18949_) );
	OAI21X1 OAI21X1_3654 ( .gnd(gnd), .vdd(vdd), .A(_18948_), .B(_17412__bF_buf1), .C(_18949_), .Y(_18950_) );
	NOR2X1 NOR2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_18947_), .B(_18950_), .Y(_18951_) );
	INVX1 INVX1_2707 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_28_), .Y(_18952_) );
	NAND3X1 NAND3X1_3712 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf1), .B(registers_r31_28_), .C(_17419__bF_buf1), .Y(_18953_) );
	OAI21X1 OAI21X1_3655 ( .gnd(gnd), .vdd(vdd), .A(_18952_), .B(_17418__bF_buf1), .C(_18953_), .Y(_18954_) );
	INVX1 INVX1_2708 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_28_), .Y(_18955_) );
	NAND3X1 NAND3X1_3713 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_28_), .B(_17392__bF_buf2), .C(_17413__bF_buf6), .Y(_18956_) );
	OAI21X1 OAI21X1_3656 ( .gnd(gnd), .vdd(vdd), .A(_18955_), .B(_17423__bF_buf1), .C(_18956_), .Y(_18957_) );
	NOR2X1 NOR2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_18954_), .B(_18957_), .Y(_18958_) );
	NAND2X1 NAND2X1_3518 ( .gnd(gnd), .vdd(vdd), .A(_18958_), .B(_18951_), .Y(_18959_) );
	NOR2X1 NOR2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_18959_), .B(_18944_), .Y(_18960_) );
	AOI22X1 AOI22X1_434 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf1), .B(registers_a2_28_), .C(registers_r1_28_), .D(_17431__bF_buf1), .Y(_18961_) );
	AOI22X1 AOI22X1_435 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf1), .B(registers_r4_28_), .C(registers_r5_28_), .D(_17436__bF_buf1), .Y(_18962_) );
	INVX1 INVX1_2709 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_28_), .Y(_18963_) );
	NAND3X1 NAND3X1_3714 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_28_), .B(_17432__bF_buf4), .C(_17392__bF_buf1), .Y(_18964_) );
	OAI21X1 OAI21X1_3657 ( .gnd(gnd), .vdd(vdd), .A(_18963_), .B(_17443__bF_buf1), .C(_18964_), .Y(_18965_) );
	AOI21X1 AOI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_28_), .B(_17440__bF_buf1), .C(_18965_), .Y(_18966_) );
	NAND3X1 NAND3X1_3715 ( .gnd(gnd), .vdd(vdd), .A(_18961_), .B(_18962_), .C(_18966_), .Y(_18967_) );
	INVX1 INVX1_2710 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_28_), .Y(_18968_) );
	INVX1 INVX1_2711 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_28_), .Y(_18969_) );
	OAI22X1 OAI22X1_380 ( .gnd(gnd), .vdd(vdd), .A(_18969_), .B(_17450__bF_buf1), .C(_18968_), .D(_17449__bF_buf1), .Y(_18970_) );
	INVX1 INVX1_2712 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_28_), .Y(_18971_) );
	INVX1 INVX1_2713 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_28_), .Y(_18972_) );
	OAI22X1 OAI22X1_381 ( .gnd(gnd), .vdd(vdd), .A(_18971_), .B(_17456__bF_buf1), .C(_18972_), .D(_17454__bF_buf1), .Y(_18973_) );
	NOR2X1 NOR2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_18973_), .B(_18970_), .Y(_18974_) );
	INVX1 INVX1_2714 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_28_), .Y(_18975_) );
	INVX1 INVX1_2715 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_28_), .Y(_18976_) );
	OAI22X1 OAI22X1_382 ( .gnd(gnd), .vdd(vdd), .A(_18975_), .B(_17461__bF_buf1), .C(_18976_), .D(_17462__bF_buf1), .Y(_18977_) );
	INVX1 INVX1_2716 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_28_), .Y(_18978_) );
	INVX1 INVX1_2717 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_28_), .Y(_18979_) );
	OAI22X1 OAI22X1_383 ( .gnd(gnd), .vdd(vdd), .A(_18979_), .B(_17467__bF_buf1), .C(_18978_), .D(_17466__bF_buf1), .Y(_18980_) );
	NOR2X1 NOR2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_18977_), .B(_18980_), .Y(_18981_) );
	NAND2X1 NAND2X1_3519 ( .gnd(gnd), .vdd(vdd), .A(_18974_), .B(_18981_), .Y(_18982_) );
	NOR2X1 NOR2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_18967_), .B(_18982_), .Y(_18983_) );
	NAND2X1 NAND2X1_3520 ( .gnd(gnd), .vdd(vdd), .A(_18983_), .B(_18960_), .Y(_428__28_) );
	NAND3X1 NAND3X1_3716 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_29_), .B(_17373__bF_buf0), .C(_17371__bF_buf4), .Y(_18984_) );
	NAND3X1 NAND3X1_3717 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_29_), .B(_17376__bF_buf0), .C(_17371__bF_buf3), .Y(_18985_) );
	NAND2X1 NAND2X1_3521 ( .gnd(gnd), .vdd(vdd), .A(_18984_), .B(_18985_), .Y(_18986_) );
	INVX1 INVX1_2718 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_29_), .Y(_18987_) );
	INVX1 INVX1_2719 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_29_), .Y(_18988_) );
	OAI22X1 OAI22X1_384 ( .gnd(gnd), .vdd(vdd), .A(_18987_), .B(_17384__bF_buf0), .C(_18988_), .D(_17383__bF_buf0), .Y(_18989_) );
	NOR2X1 NOR2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_18986_), .B(_18989_), .Y(_18990_) );
	INVX1 INVX1_2720 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_29_), .Y(_18991_) );
	INVX1 INVX1_2721 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_29_), .Y(_18992_) );
	OAI22X1 OAI22X1_385 ( .gnd(gnd), .vdd(vdd), .A(_18991_), .B(_17394__bF_buf0), .C(_18992_), .D(_17393__bF_buf0), .Y(_18993_) );
	INVX1 INVX1_2722 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_29_), .Y(_18994_) );
	INVX1 INVX1_2723 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_29_), .Y(_18995_) );
	OAI22X1 OAI22X1_386 ( .gnd(gnd), .vdd(vdd), .A(_18994_), .B(_17401__bF_buf0), .C(_18995_), .D(_17400__bF_buf0), .Y(_18996_) );
	NOR2X1 NOR2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_18996_), .B(_18993_), .Y(_18997_) );
	NAND2X1 NAND2X1_3522 ( .gnd(gnd), .vdd(vdd), .A(_18990_), .B(_18997_), .Y(_18998_) );
	INVX1 INVX1_2724 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_29_), .Y(_18999_) );
	INVX1 INVX1_2725 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_29_), .Y(_19000_) );
	OAI22X1 OAI22X1_387 ( .gnd(gnd), .vdd(vdd), .A(_19000_), .B(_17408__bF_buf0), .C(_18999_), .D(_17407__bF_buf0), .Y(_19001_) );
	INVX1 INVX1_2726 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_29_), .Y(_19002_) );
	NAND3X1 NAND3X1_3718 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_29_), .B(_17411__bF_buf2), .C(_17413__bF_buf5), .Y(_19003_) );
	OAI21X1 OAI21X1_3658 ( .gnd(gnd), .vdd(vdd), .A(_19002_), .B(_17412__bF_buf0), .C(_19003_), .Y(_19004_) );
	NOR2X1 NOR2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_19001_), .B(_19004_), .Y(_19005_) );
	INVX1 INVX1_2727 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_29_), .Y(_19006_) );
	NAND3X1 NAND3X1_3719 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf0), .B(registers_r31_29_), .C(_17419__bF_buf0), .Y(_19007_) );
	OAI21X1 OAI21X1_3659 ( .gnd(gnd), .vdd(vdd), .A(_19006_), .B(_17418__bF_buf0), .C(_19007_), .Y(_19008_) );
	INVX1 INVX1_2728 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_29_), .Y(_19009_) );
	NAND3X1 NAND3X1_3720 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_29_), .B(_17392__bF_buf0), .C(_17413__bF_buf4), .Y(_19010_) );
	OAI21X1 OAI21X1_3660 ( .gnd(gnd), .vdd(vdd), .A(_19009_), .B(_17423__bF_buf0), .C(_19010_), .Y(_19011_) );
	NOR2X1 NOR2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_19008_), .B(_19011_), .Y(_19012_) );
	NAND2X1 NAND2X1_3523 ( .gnd(gnd), .vdd(vdd), .A(_19012_), .B(_19005_), .Y(_19013_) );
	NOR2X1 NOR2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_19013_), .B(_18998_), .Y(_19014_) );
	AOI22X1 AOI22X1_436 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf0), .B(registers_a2_29_), .C(registers_r1_29_), .D(_17431__bF_buf0), .Y(_19015_) );
	AOI22X1 AOI22X1_437 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf0), .B(registers_r4_29_), .C(registers_r5_29_), .D(_17436__bF_buf0), .Y(_19016_) );
	INVX1 INVX1_2729 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_29_), .Y(_19017_) );
	NAND3X1 NAND3X1_3721 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_29_), .B(_17432__bF_buf3), .C(_17392__bF_buf7), .Y(_19018_) );
	OAI21X1 OAI21X1_3661 ( .gnd(gnd), .vdd(vdd), .A(_19017_), .B(_17443__bF_buf0), .C(_19018_), .Y(_19019_) );
	AOI21X1 AOI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_29_), .B(_17440__bF_buf0), .C(_19019_), .Y(_19020_) );
	NAND3X1 NAND3X1_3722 ( .gnd(gnd), .vdd(vdd), .A(_19015_), .B(_19016_), .C(_19020_), .Y(_19021_) );
	INVX1 INVX1_2730 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_29_), .Y(_19022_) );
	INVX1 INVX1_2731 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_29_), .Y(_19023_) );
	OAI22X1 OAI22X1_388 ( .gnd(gnd), .vdd(vdd), .A(_19023_), .B(_17450__bF_buf0), .C(_19022_), .D(_17449__bF_buf0), .Y(_19024_) );
	INVX1 INVX1_2732 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_29_), .Y(_19025_) );
	INVX1 INVX1_2733 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_29_), .Y(_19026_) );
	OAI22X1 OAI22X1_389 ( .gnd(gnd), .vdd(vdd), .A(_19025_), .B(_17456__bF_buf0), .C(_19026_), .D(_17454__bF_buf0), .Y(_19027_) );
	NOR2X1 NOR2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_19027_), .B(_19024_), .Y(_19028_) );
	INVX1 INVX1_2734 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_29_), .Y(_19029_) );
	INVX1 INVX1_2735 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_29_), .Y(_19030_) );
	OAI22X1 OAI22X1_390 ( .gnd(gnd), .vdd(vdd), .A(_19029_), .B(_17461__bF_buf0), .C(_19030_), .D(_17462__bF_buf0), .Y(_19031_) );
	INVX1 INVX1_2736 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_29_), .Y(_19032_) );
	INVX1 INVX1_2737 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_29_), .Y(_19033_) );
	OAI22X1 OAI22X1_391 ( .gnd(gnd), .vdd(vdd), .A(_19033_), .B(_17467__bF_buf0), .C(_19032_), .D(_17466__bF_buf0), .Y(_19034_) );
	NOR2X1 NOR2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_19031_), .B(_19034_), .Y(_19035_) );
	NAND2X1 NAND2X1_3524 ( .gnd(gnd), .vdd(vdd), .A(_19028_), .B(_19035_), .Y(_19036_) );
	NOR2X1 NOR2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_19021_), .B(_19036_), .Y(_19037_) );
	NAND2X1 NAND2X1_3525 ( .gnd(gnd), .vdd(vdd), .A(_19037_), .B(_19014_), .Y(_428__29_) );
	NAND3X1 NAND3X1_3723 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_30_), .B(_17373__bF_buf5), .C(_17371__bF_buf2), .Y(_19038_) );
	NAND3X1 NAND3X1_3724 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_30_), .B(_17376__bF_buf5), .C(_17371__bF_buf1), .Y(_19039_) );
	NAND2X1 NAND2X1_3526 ( .gnd(gnd), .vdd(vdd), .A(_19038_), .B(_19039_), .Y(_19040_) );
	INVX1 INVX1_2738 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_30_), .Y(_19041_) );
	INVX1 INVX1_2739 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_30_), .Y(_19042_) );
	OAI22X1 OAI22X1_392 ( .gnd(gnd), .vdd(vdd), .A(_19041_), .B(_17384__bF_buf4), .C(_19042_), .D(_17383__bF_buf4), .Y(_19043_) );
	NOR2X1 NOR2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_19040_), .B(_19043_), .Y(_19044_) );
	INVX1 INVX1_2740 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_30_), .Y(_19045_) );
	INVX1 INVX1_2741 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_30_), .Y(_19046_) );
	OAI22X1 OAI22X1_393 ( .gnd(gnd), .vdd(vdd), .A(_19045_), .B(_17394__bF_buf4), .C(_19046_), .D(_17393__bF_buf4), .Y(_19047_) );
	INVX1 INVX1_2742 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_30_), .Y(_19048_) );
	INVX1 INVX1_2743 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_30_), .Y(_19049_) );
	OAI22X1 OAI22X1_394 ( .gnd(gnd), .vdd(vdd), .A(_19048_), .B(_17401__bF_buf4), .C(_19049_), .D(_17400__bF_buf4), .Y(_19050_) );
	NOR2X1 NOR2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_19050_), .B(_19047_), .Y(_19051_) );
	NAND2X1 NAND2X1_3527 ( .gnd(gnd), .vdd(vdd), .A(_19044_), .B(_19051_), .Y(_19052_) );
	INVX1 INVX1_2744 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_30_), .Y(_19053_) );
	INVX1 INVX1_2745 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_30_), .Y(_19054_) );
	OAI22X1 OAI22X1_395 ( .gnd(gnd), .vdd(vdd), .A(_19054_), .B(_17408__bF_buf4), .C(_19053_), .D(_17407__bF_buf4), .Y(_19055_) );
	INVX1 INVX1_2746 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_30_), .Y(_19056_) );
	NAND3X1 NAND3X1_3725 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_30_), .B(_17411__bF_buf1), .C(_17413__bF_buf3), .Y(_19057_) );
	OAI21X1 OAI21X1_3662 ( .gnd(gnd), .vdd(vdd), .A(_19056_), .B(_17412__bF_buf4), .C(_19057_), .Y(_19058_) );
	NOR2X1 NOR2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_19055_), .B(_19058_), .Y(_19059_) );
	INVX1 INVX1_2747 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_30_), .Y(_19060_) );
	NAND3X1 NAND3X1_3726 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf6), .B(registers_r31_30_), .C(_17419__bF_buf4), .Y(_19061_) );
	OAI21X1 OAI21X1_3663 ( .gnd(gnd), .vdd(vdd), .A(_19060_), .B(_17418__bF_buf4), .C(_19061_), .Y(_19062_) );
	INVX1 INVX1_2748 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_30_), .Y(_19063_) );
	NAND3X1 NAND3X1_3727 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_30_), .B(_17392__bF_buf6), .C(_17413__bF_buf2), .Y(_19064_) );
	OAI21X1 OAI21X1_3664 ( .gnd(gnd), .vdd(vdd), .A(_19063_), .B(_17423__bF_buf4), .C(_19064_), .Y(_19065_) );
	NOR2X1 NOR2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_19062_), .B(_19065_), .Y(_19066_) );
	NAND2X1 NAND2X1_3528 ( .gnd(gnd), .vdd(vdd), .A(_19066_), .B(_19059_), .Y(_19067_) );
	NOR2X1 NOR2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_19067_), .B(_19052_), .Y(_19068_) );
	AOI22X1 AOI22X1_438 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf4), .B(registers_a2_30_), .C(registers_r1_30_), .D(_17431__bF_buf4), .Y(_19069_) );
	AOI22X1 AOI22X1_439 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf4), .B(registers_r4_30_), .C(registers_r5_30_), .D(_17436__bF_buf4), .Y(_19070_) );
	INVX1 INVX1_2749 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_30_), .Y(_19071_) );
	NAND3X1 NAND3X1_3728 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_30_), .B(_17432__bF_buf2), .C(_17392__bF_buf5), .Y(_19072_) );
	OAI21X1 OAI21X1_3665 ( .gnd(gnd), .vdd(vdd), .A(_19071_), .B(_17443__bF_buf4), .C(_19072_), .Y(_19073_) );
	AOI21X1 AOI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_30_), .B(_17440__bF_buf4), .C(_19073_), .Y(_19074_) );
	NAND3X1 NAND3X1_3729 ( .gnd(gnd), .vdd(vdd), .A(_19069_), .B(_19070_), .C(_19074_), .Y(_19075_) );
	INVX1 INVX1_2750 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_30_), .Y(_19076_) );
	INVX1 INVX1_2751 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_30_), .Y(_19077_) );
	OAI22X1 OAI22X1_396 ( .gnd(gnd), .vdd(vdd), .A(_19077_), .B(_17450__bF_buf4), .C(_19076_), .D(_17449__bF_buf4), .Y(_19078_) );
	INVX1 INVX1_2752 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_30_), .Y(_19079_) );
	INVX1 INVX1_2753 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_30_), .Y(_19080_) );
	OAI22X1 OAI22X1_397 ( .gnd(gnd), .vdd(vdd), .A(_19079_), .B(_17456__bF_buf4), .C(_19080_), .D(_17454__bF_buf4), .Y(_19081_) );
	NOR2X1 NOR2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_19081_), .B(_19078_), .Y(_19082_) );
	INVX1 INVX1_2754 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_30_), .Y(_19083_) );
	INVX1 INVX1_2755 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_30_), .Y(_19084_) );
	OAI22X1 OAI22X1_398 ( .gnd(gnd), .vdd(vdd), .A(_19083_), .B(_17461__bF_buf4), .C(_19084_), .D(_17462__bF_buf4), .Y(_19085_) );
	INVX1 INVX1_2756 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_30_), .Y(_19086_) );
	INVX1 INVX1_2757 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_30_), .Y(_19087_) );
	OAI22X1 OAI22X1_399 ( .gnd(gnd), .vdd(vdd), .A(_19087_), .B(_17467__bF_buf4), .C(_19086_), .D(_17466__bF_buf4), .Y(_19088_) );
	NOR2X1 NOR2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_19085_), .B(_19088_), .Y(_19089_) );
	NAND2X1 NAND2X1_3529 ( .gnd(gnd), .vdd(vdd), .A(_19082_), .B(_19089_), .Y(_19090_) );
	NOR2X1 NOR2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_19075_), .B(_19090_), .Y(_19091_) );
	NAND2X1 NAND2X1_3530 ( .gnd(gnd), .vdd(vdd), .A(_19091_), .B(_19068_), .Y(_428__30_) );
	NAND3X1 NAND3X1_3730 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_31_), .B(_17373__bF_buf4), .C(_17371__bF_buf0), .Y(_19092_) );
	NAND3X1 NAND3X1_3731 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_31_), .B(_17376__bF_buf4), .C(_17371__bF_buf7), .Y(_19093_) );
	NAND2X1 NAND2X1_3531 ( .gnd(gnd), .vdd(vdd), .A(_19092_), .B(_19093_), .Y(_19094_) );
	INVX1 INVX1_2758 ( .gnd(gnd), .vdd(vdd), .A(registers_gp_31_), .Y(_19095_) );
	INVX1 INVX1_2759 ( .gnd(gnd), .vdd(vdd), .A(registers_r2_31_), .Y(_19096_) );
	OAI22X1 OAI22X1_400 ( .gnd(gnd), .vdd(vdd), .A(_19095_), .B(_17384__bF_buf3), .C(_19096_), .D(_17383__bF_buf3), .Y(_19097_) );
	NOR2X1 NOR2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_19094_), .B(_19097_), .Y(_19098_) );
	INVX1 INVX1_2760 ( .gnd(gnd), .vdd(vdd), .A(registers_a1_31_), .Y(_19099_) );
	INVX1 INVX1_2761 ( .gnd(gnd), .vdd(vdd), .A(registers_r9_31_), .Y(_19100_) );
	OAI22X1 OAI22X1_401 ( .gnd(gnd), .vdd(vdd), .A(_19099_), .B(_17394__bF_buf3), .C(_19100_), .D(_17393__bF_buf3), .Y(_19101_) );
	INVX1 INVX1_2762 ( .gnd(gnd), .vdd(vdd), .A(registers_a4_31_), .Y(_19102_) );
	INVX1 INVX1_2763 ( .gnd(gnd), .vdd(vdd), .A(registers_a3_31_), .Y(_19103_) );
	OAI22X1 OAI22X1_402 ( .gnd(gnd), .vdd(vdd), .A(_19102_), .B(_17401__bF_buf3), .C(_19103_), .D(_17400__bF_buf3), .Y(_19104_) );
	NOR2X1 NOR2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_19104_), .B(_19101_), .Y(_19105_) );
	NAND2X1 NAND2X1_3532 ( .gnd(gnd), .vdd(vdd), .A(_19098_), .B(_19105_), .Y(_19106_) );
	INVX1 INVX1_2764 ( .gnd(gnd), .vdd(vdd), .A(registers_r18_31_), .Y(_19107_) );
	INVX1 INVX1_2765 ( .gnd(gnd), .vdd(vdd), .A(registers_r19_31_), .Y(_19108_) );
	OAI22X1 OAI22X1_403 ( .gnd(gnd), .vdd(vdd), .A(_19108_), .B(_17408__bF_buf3), .C(_19107_), .D(_17407__bF_buf3), .Y(_19109_) );
	INVX1 INVX1_2766 ( .gnd(gnd), .vdd(vdd), .A(registers_r21_31_), .Y(_19110_) );
	NAND3X1 NAND3X1_3732 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_31_), .B(_17411__bF_buf0), .C(_17413__bF_buf1), .Y(_19111_) );
	OAI21X1 OAI21X1_3666 ( .gnd(gnd), .vdd(vdd), .A(_19110_), .B(_17412__bF_buf3), .C(_19111_), .Y(_19112_) );
	NOR2X1 NOR2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_19109_), .B(_19112_), .Y(_19113_) );
	INVX1 INVX1_2767 ( .gnd(gnd), .vdd(vdd), .A(registers_r30_31_), .Y(_19114_) );
	NAND3X1 NAND3X1_3733 ( .gnd(gnd), .vdd(vdd), .A(aLoc_frameOut_4_bF_buf5), .B(registers_r31_31_), .C(_17419__bF_buf3), .Y(_19115_) );
	OAI21X1 OAI21X1_3667 ( .gnd(gnd), .vdd(vdd), .A(_19114_), .B(_17418__bF_buf3), .C(_19115_), .Y(_19116_) );
	INVX1 INVX1_2768 ( .gnd(gnd), .vdd(vdd), .A(registers_r25_31_), .Y(_19117_) );
	NAND3X1 NAND3X1_3734 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_31_), .B(_17392__bF_buf4), .C(_17413__bF_buf0), .Y(_19118_) );
	OAI21X1 OAI21X1_3668 ( .gnd(gnd), .vdd(vdd), .A(_19117_), .B(_17423__bF_buf3), .C(_19118_), .Y(_19119_) );
	NOR2X1 NOR2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_19116_), .B(_19119_), .Y(_19120_) );
	NAND2X1 NAND2X1_3533 ( .gnd(gnd), .vdd(vdd), .A(_19120_), .B(_19113_), .Y(_19121_) );
	NOR2X1 NOR2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_19121_), .B(_19106_), .Y(_19122_) );
	AOI22X1 AOI22X1_440 ( .gnd(gnd), .vdd(vdd), .A(_17433__bF_buf3), .B(registers_a2_31_), .C(registers_r1_31_), .D(_17431__bF_buf3), .Y(_19123_) );
	AOI22X1 AOI22X1_441 ( .gnd(gnd), .vdd(vdd), .A(_17435__bF_buf3), .B(registers_r4_31_), .C(registers_r5_31_), .D(_17436__bF_buf3), .Y(_19124_) );
	INVX1 INVX1_2769 ( .gnd(gnd), .vdd(vdd), .A(registers_a5_31_), .Y(_19125_) );
	NAND3X1 NAND3X1_3735 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_31_), .B(_17432__bF_buf1), .C(_17392__bF_buf3), .Y(_19126_) );
	OAI21X1 OAI21X1_3669 ( .gnd(gnd), .vdd(vdd), .A(_19125_), .B(_17443__bF_buf3), .C(_19126_), .Y(_19127_) );
	AOI21X1 AOI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_31_), .B(_17440__bF_buf3), .C(_19127_), .Y(_19128_) );
	NAND3X1 NAND3X1_3736 ( .gnd(gnd), .vdd(vdd), .A(_19123_), .B(_19124_), .C(_19128_), .Y(_19129_) );
	INVX1 INVX1_2770 ( .gnd(gnd), .vdd(vdd), .A(registers_r22_31_), .Y(_19130_) );
	INVX1 INVX1_2771 ( .gnd(gnd), .vdd(vdd), .A(registers_r23_31_), .Y(_19131_) );
	OAI22X1 OAI22X1_404 ( .gnd(gnd), .vdd(vdd), .A(_19131_), .B(_17450__bF_buf3), .C(_19130_), .D(_17449__bF_buf3), .Y(_19132_) );
	INVX1 INVX1_2772 ( .gnd(gnd), .vdd(vdd), .A(registers_a6_31_), .Y(_19133_) );
	INVX1 INVX1_2773 ( .gnd(gnd), .vdd(vdd), .A(registers_a7_31_), .Y(_19134_) );
	OAI22X1 OAI22X1_405 ( .gnd(gnd), .vdd(vdd), .A(_19133_), .B(_17456__bF_buf3), .C(_19134_), .D(_17454__bF_buf3), .Y(_19135_) );
	NOR2X1 NOR2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_19135_), .B(_19132_), .Y(_19136_) );
	INVX1 INVX1_2774 ( .gnd(gnd), .vdd(vdd), .A(registers_r28_31_), .Y(_19137_) );
	INVX1 INVX1_2775 ( .gnd(gnd), .vdd(vdd), .A(registers_r29_31_), .Y(_19138_) );
	OAI22X1 OAI22X1_406 ( .gnd(gnd), .vdd(vdd), .A(_19137_), .B(_17461__bF_buf3), .C(_19138_), .D(_17462__bF_buf3), .Y(_19139_) );
	INVX1 INVX1_2776 ( .gnd(gnd), .vdd(vdd), .A(registers_r26_31_), .Y(_19140_) );
	INVX1 INVX1_2777 ( .gnd(gnd), .vdd(vdd), .A(registers_r27_31_), .Y(_19141_) );
	OAI22X1 OAI22X1_407 ( .gnd(gnd), .vdd(vdd), .A(_19141_), .B(_17467__bF_buf3), .C(_19140_), .D(_17466__bF_buf3), .Y(_19142_) );
	NOR2X1 NOR2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_19139_), .B(_19142_), .Y(_19143_) );
	NAND2X1 NAND2X1_3534 ( .gnd(gnd), .vdd(vdd), .A(_19136_), .B(_19143_), .Y(_19144_) );
	NOR2X1 NOR2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_19129_), .B(_19144_), .Y(_19145_) );
	NAND2X1 NAND2X1_3535 ( .gnd(gnd), .vdd(vdd), .A(_19145_), .B(_19122_), .Y(_428__31_) );
	INVX1 INVX1_2778 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_0_), .Y(_19146_) );
	NAND2X1 NAND2X1_3536 ( .gnd(gnd), .vdd(vdd), .A(registers_writeEnable), .B(instructionFrame_writeSelect_out_4_), .Y(_19147_) );
	INVX4 INVX4_25 ( .gnd(gnd), .vdd(vdd), .A(_19147_), .Y(_19148_) );
	NAND2X1 NAND2X1_3537 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_3_), .B(instructionFrame_writeSelect_out_2_), .Y(_19149_) );
	NAND2X1 NAND2X1_3538 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_1_), .B(instructionFrame_writeSelect_out_0_), .Y(_19150_) );
	NOR2X1 NOR2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_19149_), .B(_19150_), .Y(_19151_) );
	NAND2X1 NAND2X1_3539 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19151_), .Y(_19152_) );
	INVX8 INVX8_73 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf10), .Y(_19153_) );
	OAI21X1 OAI21X1_3670 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf98), .Y(_19154_) );
	AOI21X1 AOI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_19146_), .B(_19152__bF_buf6), .C(_19154_), .Y(_17362__0_) );
	INVX1 INVX1_2779 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_1_), .Y(_19155_) );
	OAI21X1 OAI21X1_3671 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf97), .Y(_19156_) );
	AOI21X1 AOI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_19155_), .B(_19152__bF_buf4), .C(_19156_), .Y(_17362__1_) );
	INVX1 INVX1_2780 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_2_), .Y(_19157_) );
	OAI21X1 OAI21X1_3672 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf96), .Y(_19158_) );
	AOI21X1 AOI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_19157_), .B(_19152__bF_buf2), .C(_19158_), .Y(_17362__2_) );
	INVX1 INVX1_2781 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_3_), .Y(_19159_) );
	OAI21X1 OAI21X1_3673 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf95), .Y(_19160_) );
	AOI21X1 AOI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_19159_), .B(_19152__bF_buf0), .C(_19160_), .Y(_17362__3_) );
	INVX1 INVX1_2782 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_4_), .Y(_19161_) );
	OAI21X1 OAI21X1_3674 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf94), .Y(_19162_) );
	AOI21X1 AOI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_19161_), .B(_19152__bF_buf6), .C(_19162_), .Y(_17362__4_) );
	INVX1 INVX1_2783 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_5_), .Y(_19163_) );
	OAI21X1 OAI21X1_3675 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf93), .Y(_19164_) );
	AOI21X1 AOI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_19163_), .B(_19152__bF_buf4), .C(_19164_), .Y(_17362__5_) );
	INVX1 INVX1_2784 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_6_), .Y(_19165_) );
	OAI21X1 OAI21X1_3676 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf92), .Y(_19166_) );
	AOI21X1 AOI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_19165_), .B(_19152__bF_buf2), .C(_19166_), .Y(_17362__6_) );
	INVX1 INVX1_2785 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_7_), .Y(_19167_) );
	OAI21X1 OAI21X1_3677 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf91), .Y(_19168_) );
	AOI21X1 AOI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_19167_), .B(_19152__bF_buf0), .C(_19168_), .Y(_17362__7_) );
	INVX1 INVX1_2786 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_8_), .Y(_19169_) );
	OAI21X1 OAI21X1_3678 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf90), .Y(_19170_) );
	AOI21X1 AOI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_19169_), .B(_19152__bF_buf6), .C(_19170_), .Y(_17362__8_) );
	INVX1 INVX1_2787 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_9_), .Y(_19171_) );
	OAI21X1 OAI21X1_3679 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf89), .Y(_19172_) );
	AOI21X1 AOI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_19171_), .B(_19152__bF_buf4), .C(_19172_), .Y(_17362__9_) );
	INVX1 INVX1_2788 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_10_), .Y(_19173_) );
	OAI21X1 OAI21X1_3680 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf88), .Y(_19174_) );
	AOI21X1 AOI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_19173_), .B(_19152__bF_buf2), .C(_19174_), .Y(_17362__10_) );
	INVX1 INVX1_2789 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_11_), .Y(_19175_) );
	OAI21X1 OAI21X1_3681 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf87), .Y(_19176_) );
	AOI21X1 AOI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_19175_), .B(_19152__bF_buf0), .C(_19176_), .Y(_17362__11_) );
	INVX1 INVX1_2790 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_12_), .Y(_19177_) );
	OAI21X1 OAI21X1_3682 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf86), .Y(_19178_) );
	AOI21X1 AOI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_19177_), .B(_19152__bF_buf6), .C(_19178_), .Y(_17362__12_) );
	INVX1 INVX1_2791 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_13_), .Y(_19179_) );
	OAI21X1 OAI21X1_3683 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf85), .Y(_19180_) );
	AOI21X1 AOI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_19179_), .B(_19152__bF_buf4), .C(_19180_), .Y(_17362__13_) );
	INVX1 INVX1_2792 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_14_), .Y(_19181_) );
	OAI21X1 OAI21X1_3684 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf84), .Y(_19182_) );
	AOI21X1 AOI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_19181_), .B(_19152__bF_buf2), .C(_19182_), .Y(_17362__14_) );
	INVX1 INVX1_2793 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_15_), .Y(_19183_) );
	OAI21X1 OAI21X1_3685 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf83), .Y(_19184_) );
	AOI21X1 AOI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_19183_), .B(_19152__bF_buf0), .C(_19184_), .Y(_17362__15_) );
	INVX1 INVX1_2794 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_16_), .Y(_19185_) );
	OAI21X1 OAI21X1_3686 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf82), .Y(_19186_) );
	AOI21X1 AOI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_19185_), .B(_19152__bF_buf6), .C(_19186_), .Y(_17362__16_) );
	INVX1 INVX1_2795 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_17_), .Y(_19187_) );
	OAI21X1 OAI21X1_3687 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf81), .Y(_19188_) );
	AOI21X1 AOI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_19187_), .B(_19152__bF_buf4), .C(_19188_), .Y(_17362__17_) );
	INVX1 INVX1_2796 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_18_), .Y(_19189_) );
	OAI21X1 OAI21X1_3688 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf80), .Y(_19190_) );
	AOI21X1 AOI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_19189_), .B(_19152__bF_buf2), .C(_19190_), .Y(_17362__18_) );
	INVX1 INVX1_2797 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_19_), .Y(_19191_) );
	OAI21X1 OAI21X1_3689 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf79), .Y(_19192_) );
	AOI21X1 AOI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_19191_), .B(_19152__bF_buf0), .C(_19192_), .Y(_17362__19_) );
	INVX1 INVX1_2798 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_20_), .Y(_19193_) );
	OAI21X1 OAI21X1_3690 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf78), .Y(_19194_) );
	AOI21X1 AOI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_19193_), .B(_19152__bF_buf6), .C(_19194_), .Y(_17362__20_) );
	INVX1 INVX1_2799 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_21_), .Y(_19195_) );
	OAI21X1 OAI21X1_3691 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf77), .Y(_19196_) );
	AOI21X1 AOI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_19195_), .B(_19152__bF_buf4), .C(_19196_), .Y(_17362__21_) );
	INVX1 INVX1_2800 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_22_), .Y(_19197_) );
	OAI21X1 OAI21X1_3692 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf76), .Y(_19198_) );
	AOI21X1 AOI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_19197_), .B(_19152__bF_buf2), .C(_19198_), .Y(_17362__22_) );
	INVX1 INVX1_2801 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_23_), .Y(_19199_) );
	OAI21X1 OAI21X1_3693 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf75), .Y(_19200_) );
	AOI21X1 AOI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_19199_), .B(_19152__bF_buf0), .C(_19200_), .Y(_17362__23_) );
	INVX1 INVX1_2802 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_24_), .Y(_19201_) );
	OAI21X1 OAI21X1_3694 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf74), .Y(_19202_) );
	AOI21X1 AOI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_19201_), .B(_19152__bF_buf6), .C(_19202_), .Y(_17362__24_) );
	INVX1 INVX1_2803 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_25_), .Y(_19203_) );
	OAI21X1 OAI21X1_3695 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf73), .Y(_19204_) );
	AOI21X1 AOI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_19203_), .B(_19152__bF_buf4), .C(_19204_), .Y(_17362__25_) );
	INVX1 INVX1_2804 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_26_), .Y(_19205_) );
	OAI21X1 OAI21X1_3696 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf72), .Y(_19206_) );
	AOI21X1 AOI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_19205_), .B(_19152__bF_buf2), .C(_19206_), .Y(_17362__26_) );
	INVX1 INVX1_2805 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_27_), .Y(_19207_) );
	OAI21X1 OAI21X1_3697 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf71), .Y(_19208_) );
	AOI21X1 AOI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_19207_), .B(_19152__bF_buf0), .C(_19208_), .Y(_17362__27_) );
	INVX1 INVX1_2806 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_28_), .Y(_19209_) );
	OAI21X1 OAI21X1_3698 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_19152__bF_buf7), .C(_19153__bF_buf70), .Y(_19210_) );
	AOI21X1 AOI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_19209_), .B(_19152__bF_buf6), .C(_19210_), .Y(_17362__28_) );
	INVX1 INVX1_2807 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_29_), .Y(_19211_) );
	OAI21X1 OAI21X1_3699 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_19152__bF_buf5), .C(_19153__bF_buf69), .Y(_19212_) );
	AOI21X1 AOI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_19211_), .B(_19152__bF_buf4), .C(_19212_), .Y(_17362__29_) );
	INVX1 INVX1_2808 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_30_), .Y(_19213_) );
	OAI21X1 OAI21X1_3700 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_19152__bF_buf3), .C(_19153__bF_buf68), .Y(_19214_) );
	AOI21X1 AOI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_19213_), .B(_19152__bF_buf2), .C(_19214_), .Y(_17362__30_) );
	INVX1 INVX1_2809 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_31_), .Y(_19215_) );
	OAI21X1 OAI21X1_3701 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_19152__bF_buf1), .C(_19153__bF_buf67), .Y(_19216_) );
	AOI21X1 AOI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_19215_), .B(_19152__bF_buf0), .C(_19216_), .Y(_17362__31_) );
	INVX1 INVX1_2810 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_0_), .Y(_19217_) );
	NAND2X1 NAND2X1_3540 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_1_), .B(_19217_), .Y(_19218_) );
	NOR2X1 NOR2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_19149_), .B(_19218_), .Y(_19219_) );
	NAND2X1 NAND2X1_3541 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19219_), .Y(_19220_) );
	OAI21X1 OAI21X1_3702 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf66), .Y(_19221_) );
	AOI21X1 AOI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_17417_), .B(_19220__bF_buf6), .C(_19221_), .Y(_17361__0_) );
	OAI21X1 OAI21X1_3703 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf65), .Y(_19222_) );
	AOI21X1 AOI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_17494_), .B(_19220__bF_buf4), .C(_19222_), .Y(_17361__1_) );
	OAI21X1 OAI21X1_3704 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf64), .Y(_19223_) );
	AOI21X1 AOI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_17548_), .B(_19220__bF_buf2), .C(_19223_), .Y(_17361__2_) );
	OAI21X1 OAI21X1_3705 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf63), .Y(_19224_) );
	AOI21X1 AOI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_17602_), .B(_19220__bF_buf0), .C(_19224_), .Y(_17361__3_) );
	OAI21X1 OAI21X1_3706 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf62), .Y(_19225_) );
	AOI21X1 AOI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_17656_), .B(_19220__bF_buf6), .C(_19225_), .Y(_17361__4_) );
	OAI21X1 OAI21X1_3707 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf61), .Y(_19226_) );
	AOI21X1 AOI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_17710_), .B(_19220__bF_buf4), .C(_19226_), .Y(_17361__5_) );
	OAI21X1 OAI21X1_3708 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf60), .Y(_19227_) );
	AOI21X1 AOI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_17764_), .B(_19220__bF_buf2), .C(_19227_), .Y(_17361__6_) );
	OAI21X1 OAI21X1_3709 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf59), .Y(_19228_) );
	AOI21X1 AOI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_17818_), .B(_19220__bF_buf0), .C(_19228_), .Y(_17361__7_) );
	OAI21X1 OAI21X1_3710 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf58), .Y(_19229_) );
	AOI21X1 AOI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_17872_), .B(_19220__bF_buf6), .C(_19229_), .Y(_17361__8_) );
	OAI21X1 OAI21X1_3711 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf57), .Y(_19230_) );
	AOI21X1 AOI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_17926_), .B(_19220__bF_buf4), .C(_19230_), .Y(_17361__9_) );
	OAI21X1 OAI21X1_3712 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf56), .Y(_19231_) );
	AOI21X1 AOI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_17980_), .B(_19220__bF_buf2), .C(_19231_), .Y(_17361__10_) );
	OAI21X1 OAI21X1_3713 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf55), .Y(_19232_) );
	AOI21X1 AOI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_18034_), .B(_19220__bF_buf0), .C(_19232_), .Y(_17361__11_) );
	OAI21X1 OAI21X1_3714 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf54), .Y(_19233_) );
	AOI21X1 AOI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_18088_), .B(_19220__bF_buf6), .C(_19233_), .Y(_17361__12_) );
	OAI21X1 OAI21X1_3715 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf53), .Y(_19234_) );
	AOI21X1 AOI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_18142_), .B(_19220__bF_buf4), .C(_19234_), .Y(_17361__13_) );
	OAI21X1 OAI21X1_3716 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf52), .Y(_19235_) );
	AOI21X1 AOI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_18196_), .B(_19220__bF_buf2), .C(_19235_), .Y(_17361__14_) );
	OAI21X1 OAI21X1_3717 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf51), .Y(_19236_) );
	AOI21X1 AOI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_18250_), .B(_19220__bF_buf0), .C(_19236_), .Y(_17361__15_) );
	OAI21X1 OAI21X1_3718 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf50), .Y(_19237_) );
	AOI21X1 AOI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_18304_), .B(_19220__bF_buf6), .C(_19237_), .Y(_17361__16_) );
	OAI21X1 OAI21X1_3719 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf49), .Y(_19238_) );
	AOI21X1 AOI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_18358_), .B(_19220__bF_buf4), .C(_19238_), .Y(_17361__17_) );
	OAI21X1 OAI21X1_3720 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf48), .Y(_19239_) );
	AOI21X1 AOI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_18412_), .B(_19220__bF_buf2), .C(_19239_), .Y(_17361__18_) );
	OAI21X1 OAI21X1_3721 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf47), .Y(_19240_) );
	AOI21X1 AOI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_18466_), .B(_19220__bF_buf0), .C(_19240_), .Y(_17361__19_) );
	OAI21X1 OAI21X1_3722 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf46), .Y(_19241_) );
	AOI21X1 AOI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_18520_), .B(_19220__bF_buf6), .C(_19241_), .Y(_17361__20_) );
	OAI21X1 OAI21X1_3723 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf45), .Y(_19242_) );
	AOI21X1 AOI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_18574_), .B(_19220__bF_buf4), .C(_19242_), .Y(_17361__21_) );
	OAI21X1 OAI21X1_3724 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf44), .Y(_19243_) );
	AOI21X1 AOI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_18628_), .B(_19220__bF_buf2), .C(_19243_), .Y(_17361__22_) );
	OAI21X1 OAI21X1_3725 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf43), .Y(_19244_) );
	AOI21X1 AOI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_18682_), .B(_19220__bF_buf0), .C(_19244_), .Y(_17361__23_) );
	OAI21X1 OAI21X1_3726 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf42), .Y(_19245_) );
	AOI21X1 AOI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_18736_), .B(_19220__bF_buf6), .C(_19245_), .Y(_17361__24_) );
	OAI21X1 OAI21X1_3727 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf41), .Y(_19246_) );
	AOI21X1 AOI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_18790_), .B(_19220__bF_buf4), .C(_19246_), .Y(_17361__25_) );
	OAI21X1 OAI21X1_3728 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf40), .Y(_19247_) );
	AOI21X1 AOI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_18844_), .B(_19220__bF_buf2), .C(_19247_), .Y(_17361__26_) );
	OAI21X1 OAI21X1_3729 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf39), .Y(_19248_) );
	AOI21X1 AOI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_18898_), .B(_19220__bF_buf0), .C(_19248_), .Y(_17361__27_) );
	OAI21X1 OAI21X1_3730 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf3), .B(_19220__bF_buf7), .C(_19153__bF_buf38), .Y(_19249_) );
	AOI21X1 AOI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_18952_), .B(_19220__bF_buf6), .C(_19249_), .Y(_17361__28_) );
	OAI21X1 OAI21X1_3731 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf3), .B(_19220__bF_buf5), .C(_19153__bF_buf37), .Y(_19250_) );
	AOI21X1 AOI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_19006_), .B(_19220__bF_buf4), .C(_19250_), .Y(_17361__29_) );
	OAI21X1 OAI21X1_3732 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf3), .B(_19220__bF_buf3), .C(_19153__bF_buf36), .Y(_19251_) );
	AOI21X1 AOI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_19060_), .B(_19220__bF_buf2), .C(_19251_), .Y(_17361__30_) );
	OAI21X1 OAI21X1_3733 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf3), .B(_19220__bF_buf1), .C(_19153__bF_buf35), .Y(_19252_) );
	AOI21X1 AOI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_19114_), .B(_19220__bF_buf0), .C(_19252_), .Y(_17361__31_) );
	INVX1 INVX1_2811 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_1_), .Y(_19253_) );
	NAND2X1 NAND2X1_3542 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_0_), .B(_19253_), .Y(_19254_) );
	NOR2X1 NOR2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_19149_), .B(_19254_), .Y(_19255_) );
	NAND2X1 NAND2X1_3543 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19255_), .Y(_19256_) );
	OAI21X1 OAI21X1_3734 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf34), .Y(_19257_) );
	AOI21X1 AOI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_17460_), .B(_19256__bF_buf6), .C(_19257_), .Y(_17359__0_) );
	OAI21X1 OAI21X1_3735 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf33), .Y(_19258_) );
	AOI21X1 AOI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_17518_), .B(_19256__bF_buf4), .C(_19258_), .Y(_17359__1_) );
	OAI21X1 OAI21X1_3736 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf32), .Y(_19259_) );
	AOI21X1 AOI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_17572_), .B(_19256__bF_buf2), .C(_19259_), .Y(_17359__2_) );
	OAI21X1 OAI21X1_3737 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf31), .Y(_19260_) );
	AOI21X1 AOI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_17626_), .B(_19256__bF_buf0), .C(_19260_), .Y(_17359__3_) );
	OAI21X1 OAI21X1_3738 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf30), .Y(_19261_) );
	AOI21X1 AOI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_17680_), .B(_19256__bF_buf6), .C(_19261_), .Y(_17359__4_) );
	OAI21X1 OAI21X1_3739 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf29), .Y(_19262_) );
	AOI21X1 AOI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_17734_), .B(_19256__bF_buf4), .C(_19262_), .Y(_17359__5_) );
	OAI21X1 OAI21X1_3740 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf28), .Y(_19263_) );
	AOI21X1 AOI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_17788_), .B(_19256__bF_buf2), .C(_19263_), .Y(_17359__6_) );
	OAI21X1 OAI21X1_3741 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf27), .Y(_19264_) );
	AOI21X1 AOI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_17842_), .B(_19256__bF_buf0), .C(_19264_), .Y(_17359__7_) );
	OAI21X1 OAI21X1_3742 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf26), .Y(_19265_) );
	AOI21X1 AOI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_17896_), .B(_19256__bF_buf6), .C(_19265_), .Y(_17359__8_) );
	OAI21X1 OAI21X1_3743 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf25), .Y(_19266_) );
	AOI21X1 AOI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_17950_), .B(_19256__bF_buf4), .C(_19266_), .Y(_17359__9_) );
	OAI21X1 OAI21X1_3744 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf24), .Y(_19267_) );
	AOI21X1 AOI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_18004_), .B(_19256__bF_buf2), .C(_19267_), .Y(_17359__10_) );
	OAI21X1 OAI21X1_3745 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf23), .Y(_19268_) );
	AOI21X1 AOI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_18058_), .B(_19256__bF_buf0), .C(_19268_), .Y(_17359__11_) );
	OAI21X1 OAI21X1_3746 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf22), .Y(_19269_) );
	AOI21X1 AOI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_18112_), .B(_19256__bF_buf6), .C(_19269_), .Y(_17359__12_) );
	OAI21X1 OAI21X1_3747 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf21), .Y(_19270_) );
	AOI21X1 AOI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_18166_), .B(_19256__bF_buf4), .C(_19270_), .Y(_17359__13_) );
	OAI21X1 OAI21X1_3748 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf20), .Y(_19271_) );
	AOI21X1 AOI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_18220_), .B(_19256__bF_buf2), .C(_19271_), .Y(_17359__14_) );
	OAI21X1 OAI21X1_3749 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf19), .Y(_19272_) );
	AOI21X1 AOI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_18274_), .B(_19256__bF_buf0), .C(_19272_), .Y(_17359__15_) );
	OAI21X1 OAI21X1_3750 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf18), .Y(_19273_) );
	AOI21X1 AOI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_18328_), .B(_19256__bF_buf6), .C(_19273_), .Y(_17359__16_) );
	OAI21X1 OAI21X1_3751 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf17), .Y(_19274_) );
	AOI21X1 AOI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_18382_), .B(_19256__bF_buf4), .C(_19274_), .Y(_17359__17_) );
	OAI21X1 OAI21X1_3752 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf16), .Y(_19275_) );
	AOI21X1 AOI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_18436_), .B(_19256__bF_buf2), .C(_19275_), .Y(_17359__18_) );
	OAI21X1 OAI21X1_3753 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf15), .Y(_19276_) );
	AOI21X1 AOI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_18490_), .B(_19256__bF_buf0), .C(_19276_), .Y(_17359__19_) );
	OAI21X1 OAI21X1_3754 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf14), .Y(_19277_) );
	AOI21X1 AOI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_18544_), .B(_19256__bF_buf6), .C(_19277_), .Y(_17359__20_) );
	OAI21X1 OAI21X1_3755 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf13), .Y(_19278_) );
	AOI21X1 AOI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_18598_), .B(_19256__bF_buf4), .C(_19278_), .Y(_17359__21_) );
	OAI21X1 OAI21X1_3756 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf12), .Y(_19279_) );
	AOI21X1 AOI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_18652_), .B(_19256__bF_buf2), .C(_19279_), .Y(_17359__22_) );
	OAI21X1 OAI21X1_3757 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf11), .Y(_19280_) );
	AOI21X1 AOI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_18706_), .B(_19256__bF_buf0), .C(_19280_), .Y(_17359__23_) );
	OAI21X1 OAI21X1_3758 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf10), .Y(_19281_) );
	AOI21X1 AOI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_18760_), .B(_19256__bF_buf6), .C(_19281_), .Y(_17359__24_) );
	OAI21X1 OAI21X1_3759 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf9), .Y(_19282_) );
	AOI21X1 AOI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_18814_), .B(_19256__bF_buf4), .C(_19282_), .Y(_17359__25_) );
	OAI21X1 OAI21X1_3760 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf8), .Y(_19283_) );
	AOI21X1 AOI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_18868_), .B(_19256__bF_buf2), .C(_19283_), .Y(_17359__26_) );
	OAI21X1 OAI21X1_3761 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf7), .Y(_19284_) );
	AOI21X1 AOI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_18922_), .B(_19256__bF_buf0), .C(_19284_), .Y(_17359__27_) );
	OAI21X1 OAI21X1_3762 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf2), .B(_19256__bF_buf7), .C(_19153__bF_buf6), .Y(_19285_) );
	AOI21X1 AOI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_18976_), .B(_19256__bF_buf6), .C(_19285_), .Y(_17359__28_) );
	OAI21X1 OAI21X1_3763 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf2), .B(_19256__bF_buf5), .C(_19153__bF_buf5), .Y(_19286_) );
	AOI21X1 AOI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_19030_), .B(_19256__bF_buf4), .C(_19286_), .Y(_17359__29_) );
	OAI21X1 OAI21X1_3764 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf2), .B(_19256__bF_buf3), .C(_19153__bF_buf4), .Y(_19287_) );
	AOI21X1 AOI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_19084_), .B(_19256__bF_buf2), .C(_19287_), .Y(_17359__30_) );
	OAI21X1 OAI21X1_3765 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf2), .B(_19256__bF_buf1), .C(_19153__bF_buf3), .Y(_19288_) );
	AOI21X1 AOI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_19138_), .B(_19256__bF_buf0), .C(_19288_), .Y(_17359__31_) );
	NOR2X1 NOR2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_1_), .B(instructionFrame_writeSelect_out_0_), .Y(_19289_) );
	INVX1 INVX1_2812 ( .gnd(gnd), .vdd(vdd), .A(_19289_), .Y(_19290_) );
	NOR2X1 NOR2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_19149_), .B(_19290_), .Y(_19291_) );
	NAND2X1 NAND2X1_3544 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19291_), .Y(_19292_) );
	OAI21X1 OAI21X1_3766 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf2), .Y(_19293_) );
	AOI21X1 AOI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_17459_), .B(_19292__bF_buf6), .C(_19293_), .Y(_17358__0_) );
	OAI21X1 OAI21X1_3767 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf1), .Y(_19294_) );
	AOI21X1 AOI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_17517_), .B(_19292__bF_buf4), .C(_19294_), .Y(_17358__1_) );
	OAI21X1 OAI21X1_3768 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf0), .Y(_19295_) );
	AOI21X1 AOI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_17571_), .B(_19292__bF_buf2), .C(_19295_), .Y(_17358__2_) );
	OAI21X1 OAI21X1_3769 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf98), .Y(_19296_) );
	AOI21X1 AOI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_17625_), .B(_19292__bF_buf0), .C(_19296_), .Y(_17358__3_) );
	OAI21X1 OAI21X1_3770 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf97), .Y(_19297_) );
	AOI21X1 AOI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_17679_), .B(_19292__bF_buf6), .C(_19297_), .Y(_17358__4_) );
	OAI21X1 OAI21X1_3771 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf96), .Y(_19298_) );
	AOI21X1 AOI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_17733_), .B(_19292__bF_buf4), .C(_19298_), .Y(_17358__5_) );
	OAI21X1 OAI21X1_3772 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf95), .Y(_19299_) );
	AOI21X1 AOI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_17787_), .B(_19292__bF_buf2), .C(_19299_), .Y(_17358__6_) );
	OAI21X1 OAI21X1_3773 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf94), .Y(_19300_) );
	AOI21X1 AOI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_17841_), .B(_19292__bF_buf0), .C(_19300_), .Y(_17358__7_) );
	OAI21X1 OAI21X1_3774 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf93), .Y(_19301_) );
	AOI21X1 AOI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_17895_), .B(_19292__bF_buf6), .C(_19301_), .Y(_17358__8_) );
	OAI21X1 OAI21X1_3775 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf92), .Y(_19302_) );
	AOI21X1 AOI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_17949_), .B(_19292__bF_buf4), .C(_19302_), .Y(_17358__9_) );
	OAI21X1 OAI21X1_3776 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf91), .Y(_19303_) );
	AOI21X1 AOI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_18003_), .B(_19292__bF_buf2), .C(_19303_), .Y(_17358__10_) );
	OAI21X1 OAI21X1_3777 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf90), .Y(_19304_) );
	AOI21X1 AOI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_18057_), .B(_19292__bF_buf0), .C(_19304_), .Y(_17358__11_) );
	OAI21X1 OAI21X1_3778 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf89), .Y(_19305_) );
	AOI21X1 AOI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_18111_), .B(_19292__bF_buf6), .C(_19305_), .Y(_17358__12_) );
	OAI21X1 OAI21X1_3779 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf88), .Y(_19306_) );
	AOI21X1 AOI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_18165_), .B(_19292__bF_buf4), .C(_19306_), .Y(_17358__13_) );
	OAI21X1 OAI21X1_3780 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf87), .Y(_19307_) );
	AOI21X1 AOI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_18219_), .B(_19292__bF_buf2), .C(_19307_), .Y(_17358__14_) );
	OAI21X1 OAI21X1_3781 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf86), .Y(_19308_) );
	AOI21X1 AOI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_18273_), .B(_19292__bF_buf0), .C(_19308_), .Y(_17358__15_) );
	OAI21X1 OAI21X1_3782 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf85), .Y(_19309_) );
	AOI21X1 AOI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_18327_), .B(_19292__bF_buf6), .C(_19309_), .Y(_17358__16_) );
	OAI21X1 OAI21X1_3783 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf84), .Y(_19310_) );
	AOI21X1 AOI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_18381_), .B(_19292__bF_buf4), .C(_19310_), .Y(_17358__17_) );
	OAI21X1 OAI21X1_3784 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf83), .Y(_19311_) );
	AOI21X1 AOI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_18435_), .B(_19292__bF_buf2), .C(_19311_), .Y(_17358__18_) );
	OAI21X1 OAI21X1_3785 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf82), .Y(_19312_) );
	AOI21X1 AOI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_18489_), .B(_19292__bF_buf0), .C(_19312_), .Y(_17358__19_) );
	OAI21X1 OAI21X1_3786 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf81), .Y(_19313_) );
	AOI21X1 AOI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_18543_), .B(_19292__bF_buf6), .C(_19313_), .Y(_17358__20_) );
	OAI21X1 OAI21X1_3787 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf80), .Y(_19314_) );
	AOI21X1 AOI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_18597_), .B(_19292__bF_buf4), .C(_19314_), .Y(_17358__21_) );
	OAI21X1 OAI21X1_3788 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf79), .Y(_19315_) );
	AOI21X1 AOI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_18651_), .B(_19292__bF_buf2), .C(_19315_), .Y(_17358__22_) );
	OAI21X1 OAI21X1_3789 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf78), .Y(_19316_) );
	AOI21X1 AOI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_18705_), .B(_19292__bF_buf0), .C(_19316_), .Y(_17358__23_) );
	OAI21X1 OAI21X1_3790 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf77), .Y(_19317_) );
	AOI21X1 AOI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_18759_), .B(_19292__bF_buf6), .C(_19317_), .Y(_17358__24_) );
	OAI21X1 OAI21X1_3791 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf76), .Y(_19318_) );
	AOI21X1 AOI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_18813_), .B(_19292__bF_buf4), .C(_19318_), .Y(_17358__25_) );
	OAI21X1 OAI21X1_3792 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf75), .Y(_19319_) );
	AOI21X1 AOI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_18867_), .B(_19292__bF_buf2), .C(_19319_), .Y(_17358__26_) );
	OAI21X1 OAI21X1_3793 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf74), .Y(_19320_) );
	AOI21X1 AOI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_18921_), .B(_19292__bF_buf0), .C(_19320_), .Y(_17358__27_) );
	OAI21X1 OAI21X1_3794 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf1), .B(_19292__bF_buf7), .C(_19153__bF_buf73), .Y(_19321_) );
	AOI21X1 AOI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_18975_), .B(_19292__bF_buf6), .C(_19321_), .Y(_17358__28_) );
	OAI21X1 OAI21X1_3795 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf1), .B(_19292__bF_buf5), .C(_19153__bF_buf72), .Y(_19322_) );
	AOI21X1 AOI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_19029_), .B(_19292__bF_buf4), .C(_19322_), .Y(_17358__29_) );
	OAI21X1 OAI21X1_3796 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf1), .B(_19292__bF_buf3), .C(_19153__bF_buf71), .Y(_19323_) );
	AOI21X1 AOI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_19083_), .B(_19292__bF_buf2), .C(_19323_), .Y(_17358__30_) );
	OAI21X1 OAI21X1_3797 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf1), .B(_19292__bF_buf1), .C(_19153__bF_buf70), .Y(_19324_) );
	AOI21X1 AOI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_19137_), .B(_19292__bF_buf0), .C(_19324_), .Y(_17358__31_) );
	INVX1 INVX1_2813 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_2_), .Y(_19325_) );
	NAND2X1 NAND2X1_3545 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_3_), .B(_19325_), .Y(_19326_) );
	NOR2X1 NOR2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_19150_), .B(_19326_), .Y(_19327_) );
	NAND2X1 NAND2X1_3546 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19327_), .Y(_19328_) );
	OAI21X1 OAI21X1_3798 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf69), .Y(_19329_) );
	AOI21X1 AOI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_17465_), .B(_19328__bF_buf6), .C(_19329_), .Y(_17357__0_) );
	OAI21X1 OAI21X1_3799 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf68), .Y(_19330_) );
	AOI21X1 AOI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_17521_), .B(_19328__bF_buf4), .C(_19330_), .Y(_17357__1_) );
	OAI21X1 OAI21X1_3800 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf67), .Y(_19331_) );
	AOI21X1 AOI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_17575_), .B(_19328__bF_buf2), .C(_19331_), .Y(_17357__2_) );
	OAI21X1 OAI21X1_3801 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf66), .Y(_19332_) );
	AOI21X1 AOI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_17629_), .B(_19328__bF_buf0), .C(_19332_), .Y(_17357__3_) );
	OAI21X1 OAI21X1_3802 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf65), .Y(_19333_) );
	AOI21X1 AOI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_17683_), .B(_19328__bF_buf6), .C(_19333_), .Y(_17357__4_) );
	OAI21X1 OAI21X1_3803 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf64), .Y(_19334_) );
	AOI21X1 AOI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_17737_), .B(_19328__bF_buf4), .C(_19334_), .Y(_17357__5_) );
	OAI21X1 OAI21X1_3804 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf63), .Y(_19335_) );
	AOI21X1 AOI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_17791_), .B(_19328__bF_buf2), .C(_19335_), .Y(_17357__6_) );
	OAI21X1 OAI21X1_3805 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf62), .Y(_19336_) );
	AOI21X1 AOI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_17845_), .B(_19328__bF_buf0), .C(_19336_), .Y(_17357__7_) );
	OAI21X1 OAI21X1_3806 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf61), .Y(_19337_) );
	AOI21X1 AOI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_17899_), .B(_19328__bF_buf6), .C(_19337_), .Y(_17357__8_) );
	OAI21X1 OAI21X1_3807 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf60), .Y(_19338_) );
	AOI21X1 AOI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_17953_), .B(_19328__bF_buf4), .C(_19338_), .Y(_17357__9_) );
	OAI21X1 OAI21X1_3808 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf59), .Y(_19339_) );
	AOI21X1 AOI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_18007_), .B(_19328__bF_buf2), .C(_19339_), .Y(_17357__10_) );
	OAI21X1 OAI21X1_3809 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf58), .Y(_19340_) );
	AOI21X1 AOI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_18061_), .B(_19328__bF_buf0), .C(_19340_), .Y(_17357__11_) );
	OAI21X1 OAI21X1_3810 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf57), .Y(_19341_) );
	AOI21X1 AOI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_18115_), .B(_19328__bF_buf6), .C(_19341_), .Y(_17357__12_) );
	OAI21X1 OAI21X1_3811 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf56), .Y(_19342_) );
	AOI21X1 AOI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_18169_), .B(_19328__bF_buf4), .C(_19342_), .Y(_17357__13_) );
	OAI21X1 OAI21X1_3812 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf55), .Y(_19343_) );
	AOI21X1 AOI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_18223_), .B(_19328__bF_buf2), .C(_19343_), .Y(_17357__14_) );
	OAI21X1 OAI21X1_3813 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf54), .Y(_19344_) );
	AOI21X1 AOI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_18277_), .B(_19328__bF_buf0), .C(_19344_), .Y(_17357__15_) );
	OAI21X1 OAI21X1_3814 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf53), .Y(_19345_) );
	AOI21X1 AOI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_18331_), .B(_19328__bF_buf6), .C(_19345_), .Y(_17357__16_) );
	OAI21X1 OAI21X1_3815 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf52), .Y(_19346_) );
	AOI21X1 AOI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_18385_), .B(_19328__bF_buf4), .C(_19346_), .Y(_17357__17_) );
	OAI21X1 OAI21X1_3816 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf51), .Y(_19347_) );
	AOI21X1 AOI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_18439_), .B(_19328__bF_buf2), .C(_19347_), .Y(_17357__18_) );
	OAI21X1 OAI21X1_3817 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf50), .Y(_19348_) );
	AOI21X1 AOI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_18493_), .B(_19328__bF_buf0), .C(_19348_), .Y(_17357__19_) );
	OAI21X1 OAI21X1_3818 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf49), .Y(_19349_) );
	AOI21X1 AOI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_18547_), .B(_19328__bF_buf6), .C(_19349_), .Y(_17357__20_) );
	OAI21X1 OAI21X1_3819 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf48), .Y(_19350_) );
	AOI21X1 AOI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_18601_), .B(_19328__bF_buf4), .C(_19350_), .Y(_17357__21_) );
	OAI21X1 OAI21X1_3820 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf47), .Y(_19351_) );
	AOI21X1 AOI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_18655_), .B(_19328__bF_buf2), .C(_19351_), .Y(_17357__22_) );
	OAI21X1 OAI21X1_3821 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf46), .Y(_19352_) );
	AOI21X1 AOI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_18709_), .B(_19328__bF_buf0), .C(_19352_), .Y(_17357__23_) );
	OAI21X1 OAI21X1_3822 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf45), .Y(_19353_) );
	AOI21X1 AOI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_18763_), .B(_19328__bF_buf6), .C(_19353_), .Y(_17357__24_) );
	OAI21X1 OAI21X1_3823 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf44), .Y(_19354_) );
	AOI21X1 AOI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_18817_), .B(_19328__bF_buf4), .C(_19354_), .Y(_17357__25_) );
	OAI21X1 OAI21X1_3824 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf43), .Y(_19355_) );
	AOI21X1 AOI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_18871_), .B(_19328__bF_buf2), .C(_19355_), .Y(_17357__26_) );
	OAI21X1 OAI21X1_3825 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf42), .Y(_19356_) );
	AOI21X1 AOI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_18925_), .B(_19328__bF_buf0), .C(_19356_), .Y(_17357__27_) );
	OAI21X1 OAI21X1_3826 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf0), .B(_19328__bF_buf7), .C(_19153__bF_buf41), .Y(_19357_) );
	AOI21X1 AOI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_18979_), .B(_19328__bF_buf6), .C(_19357_), .Y(_17357__28_) );
	OAI21X1 OAI21X1_3827 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf0), .B(_19328__bF_buf5), .C(_19153__bF_buf40), .Y(_19358_) );
	AOI21X1 AOI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_19033_), .B(_19328__bF_buf4), .C(_19358_), .Y(_17357__29_) );
	OAI21X1 OAI21X1_3828 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf0), .B(_19328__bF_buf3), .C(_19153__bF_buf39), .Y(_19359_) );
	AOI21X1 AOI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_19087_), .B(_19328__bF_buf2), .C(_19359_), .Y(_17357__30_) );
	OAI21X1 OAI21X1_3829 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf0), .B(_19328__bF_buf1), .C(_19153__bF_buf38), .Y(_19360_) );
	AOI21X1 AOI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_19141_), .B(_19328__bF_buf0), .C(_19360_), .Y(_17357__31_) );
	NOR2X1 NOR2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_19218_), .B(_19326_), .Y(_19361_) );
	NAND2X1 NAND2X1_3547 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19361_), .Y(_19362_) );
	OAI21X1 OAI21X1_3830 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf37), .Y(_19363_) );
	AOI21X1 AOI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_17464_), .B(_19362__bF_buf6), .C(_19363_), .Y(_17356__0_) );
	OAI21X1 OAI21X1_3831 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf36), .Y(_19364_) );
	AOI21X1 AOI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_17520_), .B(_19362__bF_buf4), .C(_19364_), .Y(_17356__1_) );
	OAI21X1 OAI21X1_3832 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf35), .Y(_19365_) );
	AOI21X1 AOI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_17574_), .B(_19362__bF_buf2), .C(_19365_), .Y(_17356__2_) );
	OAI21X1 OAI21X1_3833 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf34), .Y(_19366_) );
	AOI21X1 AOI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_17628_), .B(_19362__bF_buf0), .C(_19366_), .Y(_17356__3_) );
	OAI21X1 OAI21X1_3834 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf33), .Y(_19367_) );
	AOI21X1 AOI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_17682_), .B(_19362__bF_buf6), .C(_19367_), .Y(_17356__4_) );
	OAI21X1 OAI21X1_3835 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf32), .Y(_19368_) );
	AOI21X1 AOI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_17736_), .B(_19362__bF_buf4), .C(_19368_), .Y(_17356__5_) );
	OAI21X1 OAI21X1_3836 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf31), .Y(_19369_) );
	AOI21X1 AOI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_17790_), .B(_19362__bF_buf2), .C(_19369_), .Y(_17356__6_) );
	OAI21X1 OAI21X1_3837 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf30), .Y(_19370_) );
	AOI21X1 AOI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_17844_), .B(_19362__bF_buf0), .C(_19370_), .Y(_17356__7_) );
	OAI21X1 OAI21X1_3838 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf29), .Y(_19371_) );
	AOI21X1 AOI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_17898_), .B(_19362__bF_buf6), .C(_19371_), .Y(_17356__8_) );
	OAI21X1 OAI21X1_3839 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf28), .Y(_19372_) );
	AOI21X1 AOI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_17952_), .B(_19362__bF_buf4), .C(_19372_), .Y(_17356__9_) );
	OAI21X1 OAI21X1_3840 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf27), .Y(_19373_) );
	AOI21X1 AOI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_18006_), .B(_19362__bF_buf2), .C(_19373_), .Y(_17356__10_) );
	OAI21X1 OAI21X1_3841 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf26), .Y(_19374_) );
	AOI21X1 AOI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_18060_), .B(_19362__bF_buf0), .C(_19374_), .Y(_17356__11_) );
	OAI21X1 OAI21X1_3842 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf25), .Y(_19375_) );
	AOI21X1 AOI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_18114_), .B(_19362__bF_buf6), .C(_19375_), .Y(_17356__12_) );
	OAI21X1 OAI21X1_3843 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf24), .Y(_19376_) );
	AOI21X1 AOI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_18168_), .B(_19362__bF_buf4), .C(_19376_), .Y(_17356__13_) );
	OAI21X1 OAI21X1_3844 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf23), .Y(_19377_) );
	AOI21X1 AOI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_18222_), .B(_19362__bF_buf2), .C(_19377_), .Y(_17356__14_) );
	OAI21X1 OAI21X1_3845 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf22), .Y(_19378_) );
	AOI21X1 AOI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_18276_), .B(_19362__bF_buf0), .C(_19378_), .Y(_17356__15_) );
	OAI21X1 OAI21X1_3846 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf21), .Y(_19379_) );
	AOI21X1 AOI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_18330_), .B(_19362__bF_buf6), .C(_19379_), .Y(_17356__16_) );
	OAI21X1 OAI21X1_3847 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf20), .Y(_19380_) );
	AOI21X1 AOI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_18384_), .B(_19362__bF_buf4), .C(_19380_), .Y(_17356__17_) );
	OAI21X1 OAI21X1_3848 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf19), .Y(_19381_) );
	AOI21X1 AOI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_18438_), .B(_19362__bF_buf2), .C(_19381_), .Y(_17356__18_) );
	OAI21X1 OAI21X1_3849 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf18), .Y(_19382_) );
	AOI21X1 AOI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_18492_), .B(_19362__bF_buf0), .C(_19382_), .Y(_17356__19_) );
	OAI21X1 OAI21X1_3850 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf17), .Y(_19383_) );
	AOI21X1 AOI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_18546_), .B(_19362__bF_buf6), .C(_19383_), .Y(_17356__20_) );
	OAI21X1 OAI21X1_3851 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf16), .Y(_19384_) );
	AOI21X1 AOI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_18600_), .B(_19362__bF_buf4), .C(_19384_), .Y(_17356__21_) );
	OAI21X1 OAI21X1_3852 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf15), .Y(_19385_) );
	AOI21X1 AOI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_18654_), .B(_19362__bF_buf2), .C(_19385_), .Y(_17356__22_) );
	OAI21X1 OAI21X1_3853 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf14), .Y(_19386_) );
	AOI21X1 AOI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_18708_), .B(_19362__bF_buf0), .C(_19386_), .Y(_17356__23_) );
	OAI21X1 OAI21X1_3854 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf13), .Y(_19387_) );
	AOI21X1 AOI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_18762_), .B(_19362__bF_buf6), .C(_19387_), .Y(_17356__24_) );
	OAI21X1 OAI21X1_3855 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf12), .Y(_19388_) );
	AOI21X1 AOI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_18816_), .B(_19362__bF_buf4), .C(_19388_), .Y(_17356__25_) );
	OAI21X1 OAI21X1_3856 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf11), .Y(_19389_) );
	AOI21X1 AOI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_18870_), .B(_19362__bF_buf2), .C(_19389_), .Y(_17356__26_) );
	OAI21X1 OAI21X1_3857 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf10), .Y(_19390_) );
	AOI21X1 AOI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_18924_), .B(_19362__bF_buf0), .C(_19390_), .Y(_17356__27_) );
	OAI21X1 OAI21X1_3858 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_19362__bF_buf7), .C(_19153__bF_buf9), .Y(_19391_) );
	AOI21X1 AOI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_18978_), .B(_19362__bF_buf6), .C(_19391_), .Y(_17356__28_) );
	OAI21X1 OAI21X1_3859 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_19362__bF_buf5), .C(_19153__bF_buf8), .Y(_19392_) );
	AOI21X1 AOI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_19032_), .B(_19362__bF_buf4), .C(_19392_), .Y(_17356__29_) );
	OAI21X1 OAI21X1_3860 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_19362__bF_buf3), .C(_19153__bF_buf7), .Y(_19393_) );
	AOI21X1 AOI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_19086_), .B(_19362__bF_buf2), .C(_19393_), .Y(_17356__30_) );
	OAI21X1 OAI21X1_3861 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_19362__bF_buf1), .C(_19153__bF_buf6), .Y(_19394_) );
	AOI21X1 AOI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_19140_), .B(_19362__bF_buf0), .C(_19394_), .Y(_17356__31_) );
	NOR2X1 NOR2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_19254_), .B(_19326_), .Y(_19395_) );
	NAND2X1 NAND2X1_3548 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19395_), .Y(_19396_) );
	OAI21X1 OAI21X1_3862 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf5), .Y(_19397_) );
	AOI21X1 AOI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_17422_), .B(_19396__bF_buf6), .C(_19397_), .Y(_17355__0_) );
	OAI21X1 OAI21X1_3863 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf4), .Y(_19398_) );
	AOI21X1 AOI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_17497_), .B(_19396__bF_buf4), .C(_19398_), .Y(_17355__1_) );
	OAI21X1 OAI21X1_3864 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf3), .Y(_19399_) );
	AOI21X1 AOI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_17551_), .B(_19396__bF_buf2), .C(_19399_), .Y(_17355__2_) );
	OAI21X1 OAI21X1_3865 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf2), .Y(_19400_) );
	AOI21X1 AOI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_17605_), .B(_19396__bF_buf0), .C(_19400_), .Y(_17355__3_) );
	OAI21X1 OAI21X1_3866 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf1), .Y(_19401_) );
	AOI21X1 AOI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_17659_), .B(_19396__bF_buf6), .C(_19401_), .Y(_17355__4_) );
	OAI21X1 OAI21X1_3867 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf0), .Y(_19402_) );
	AOI21X1 AOI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_17713_), .B(_19396__bF_buf4), .C(_19402_), .Y(_17355__5_) );
	OAI21X1 OAI21X1_3868 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf98), .Y(_19403_) );
	AOI21X1 AOI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_17767_), .B(_19396__bF_buf2), .C(_19403_), .Y(_17355__6_) );
	OAI21X1 OAI21X1_3869 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf97), .Y(_19404_) );
	AOI21X1 AOI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_17821_), .B(_19396__bF_buf0), .C(_19404_), .Y(_17355__7_) );
	OAI21X1 OAI21X1_3870 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf96), .Y(_19405_) );
	AOI21X1 AOI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_17875_), .B(_19396__bF_buf6), .C(_19405_), .Y(_17355__8_) );
	OAI21X1 OAI21X1_3871 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf95), .Y(_19406_) );
	AOI21X1 AOI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_17929_), .B(_19396__bF_buf4), .C(_19406_), .Y(_17355__9_) );
	OAI21X1 OAI21X1_3872 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf94), .Y(_19407_) );
	AOI21X1 AOI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_17983_), .B(_19396__bF_buf2), .C(_19407_), .Y(_17355__10_) );
	OAI21X1 OAI21X1_3873 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf93), .Y(_19408_) );
	AOI21X1 AOI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_18037_), .B(_19396__bF_buf0), .C(_19408_), .Y(_17355__11_) );
	OAI21X1 OAI21X1_3874 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf92), .Y(_19409_) );
	AOI21X1 AOI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_18091_), .B(_19396__bF_buf6), .C(_19409_), .Y(_17355__12_) );
	OAI21X1 OAI21X1_3875 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf91), .Y(_19410_) );
	AOI21X1 AOI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_18145_), .B(_19396__bF_buf4), .C(_19410_), .Y(_17355__13_) );
	OAI21X1 OAI21X1_3876 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf90), .Y(_19411_) );
	AOI21X1 AOI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_18199_), .B(_19396__bF_buf2), .C(_19411_), .Y(_17355__14_) );
	OAI21X1 OAI21X1_3877 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf89), .Y(_19412_) );
	AOI21X1 AOI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_18253_), .B(_19396__bF_buf0), .C(_19412_), .Y(_17355__15_) );
	OAI21X1 OAI21X1_3878 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf88), .Y(_19413_) );
	AOI21X1 AOI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_18307_), .B(_19396__bF_buf6), .C(_19413_), .Y(_17355__16_) );
	OAI21X1 OAI21X1_3879 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf87), .Y(_19414_) );
	AOI21X1 AOI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_18361_), .B(_19396__bF_buf4), .C(_19414_), .Y(_17355__17_) );
	OAI21X1 OAI21X1_3880 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf86), .Y(_19415_) );
	AOI21X1 AOI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_18415_), .B(_19396__bF_buf2), .C(_19415_), .Y(_17355__18_) );
	OAI21X1 OAI21X1_3881 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf85), .Y(_19416_) );
	AOI21X1 AOI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_18469_), .B(_19396__bF_buf0), .C(_19416_), .Y(_17355__19_) );
	OAI21X1 OAI21X1_3882 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf84), .Y(_19417_) );
	AOI21X1 AOI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_18523_), .B(_19396__bF_buf6), .C(_19417_), .Y(_17355__20_) );
	OAI21X1 OAI21X1_3883 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf83), .Y(_19418_) );
	AOI21X1 AOI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_18577_), .B(_19396__bF_buf4), .C(_19418_), .Y(_17355__21_) );
	OAI21X1 OAI21X1_3884 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf82), .Y(_19419_) );
	AOI21X1 AOI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_18631_), .B(_19396__bF_buf2), .C(_19419_), .Y(_17355__22_) );
	OAI21X1 OAI21X1_3885 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf81), .Y(_19420_) );
	AOI21X1 AOI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_18685_), .B(_19396__bF_buf0), .C(_19420_), .Y(_17355__23_) );
	OAI21X1 OAI21X1_3886 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf80), .Y(_19421_) );
	AOI21X1 AOI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_18739_), .B(_19396__bF_buf6), .C(_19421_), .Y(_17355__24_) );
	OAI21X1 OAI21X1_3887 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf79), .Y(_19422_) );
	AOI21X1 AOI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_18793_), .B(_19396__bF_buf4), .C(_19422_), .Y(_17355__25_) );
	OAI21X1 OAI21X1_3888 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf78), .Y(_19423_) );
	AOI21X1 AOI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_18847_), .B(_19396__bF_buf2), .C(_19423_), .Y(_17355__26_) );
	OAI21X1 OAI21X1_3889 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf77), .Y(_19424_) );
	AOI21X1 AOI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_18901_), .B(_19396__bF_buf0), .C(_19424_), .Y(_17355__27_) );
	OAI21X1 OAI21X1_3890 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf3), .B(_19396__bF_buf7), .C(_19153__bF_buf76), .Y(_19425_) );
	AOI21X1 AOI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_18955_), .B(_19396__bF_buf6), .C(_19425_), .Y(_17355__28_) );
	OAI21X1 OAI21X1_3891 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf3), .B(_19396__bF_buf5), .C(_19153__bF_buf75), .Y(_19426_) );
	AOI21X1 AOI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_19009_), .B(_19396__bF_buf4), .C(_19426_), .Y(_17355__29_) );
	OAI21X1 OAI21X1_3892 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf3), .B(_19396__bF_buf3), .C(_19153__bF_buf74), .Y(_19427_) );
	AOI21X1 AOI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_19063_), .B(_19396__bF_buf2), .C(_19427_), .Y(_17355__30_) );
	OAI21X1 OAI21X1_3893 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf3), .B(_19396__bF_buf1), .C(_19153__bF_buf73), .Y(_19428_) );
	AOI21X1 AOI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_19117_), .B(_19396__bF_buf0), .C(_19428_), .Y(_17355__31_) );
	INVX1 INVX1_2814 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_0_), .Y(_19429_) );
	NOR2X1 NOR2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_19147_), .B(_19290_), .Y(_19430_) );
	INVX1 INVX1_2815 ( .gnd(gnd), .vdd(vdd), .A(_19326_), .Y(_19431_) );
	NAND2X1 NAND2X1_3549 ( .gnd(gnd), .vdd(vdd), .A(_19431_), .B(_19430_), .Y(_19432_) );
	OAI21X1 OAI21X1_3894 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf72), .Y(_19433_) );
	AOI21X1 AOI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_19429_), .B(_19432__bF_buf6), .C(_19433_), .Y(_17354__0_) );
	INVX1 INVX1_2816 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_1_), .Y(_19434_) );
	OAI21X1 OAI21X1_3895 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf71), .Y(_19435_) );
	AOI21X1 AOI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_19434_), .B(_19432__bF_buf4), .C(_19435_), .Y(_17354__1_) );
	INVX1 INVX1_2817 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_2_), .Y(_19436_) );
	OAI21X1 OAI21X1_3896 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf70), .Y(_19437_) );
	AOI21X1 AOI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_19436_), .B(_19432__bF_buf2), .C(_19437_), .Y(_17354__2_) );
	INVX1 INVX1_2818 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_3_), .Y(_19438_) );
	OAI21X1 OAI21X1_3897 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf69), .Y(_19439_) );
	AOI21X1 AOI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_19438_), .B(_19432__bF_buf0), .C(_19439_), .Y(_17354__3_) );
	INVX1 INVX1_2819 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_4_), .Y(_19440_) );
	OAI21X1 OAI21X1_3898 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf68), .Y(_19441_) );
	AOI21X1 AOI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_19440_), .B(_19432__bF_buf6), .C(_19441_), .Y(_17354__4_) );
	INVX1 INVX1_2820 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_5_), .Y(_19442_) );
	OAI21X1 OAI21X1_3899 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf67), .Y(_19443_) );
	AOI21X1 AOI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_19442_), .B(_19432__bF_buf4), .C(_19443_), .Y(_17354__5_) );
	INVX1 INVX1_2821 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_6_), .Y(_19444_) );
	OAI21X1 OAI21X1_3900 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf66), .Y(_19445_) );
	AOI21X1 AOI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_19444_), .B(_19432__bF_buf2), .C(_19445_), .Y(_17354__6_) );
	INVX1 INVX1_2822 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_7_), .Y(_19446_) );
	OAI21X1 OAI21X1_3901 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf65), .Y(_19447_) );
	AOI21X1 AOI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_19446_), .B(_19432__bF_buf0), .C(_19447_), .Y(_17354__7_) );
	INVX1 INVX1_2823 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_8_), .Y(_19448_) );
	OAI21X1 OAI21X1_3902 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf64), .Y(_19449_) );
	AOI21X1 AOI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_19448_), .B(_19432__bF_buf6), .C(_19449_), .Y(_17354__8_) );
	INVX1 INVX1_2824 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_9_), .Y(_19450_) );
	OAI21X1 OAI21X1_3903 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf63), .Y(_19451_) );
	AOI21X1 AOI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_19450_), .B(_19432__bF_buf4), .C(_19451_), .Y(_17354__9_) );
	INVX1 INVX1_2825 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_10_), .Y(_19452_) );
	OAI21X1 OAI21X1_3904 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf62), .Y(_19453_) );
	AOI21X1 AOI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_19452_), .B(_19432__bF_buf2), .C(_19453_), .Y(_17354__10_) );
	INVX1 INVX1_2826 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_11_), .Y(_19454_) );
	OAI21X1 OAI21X1_3905 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf61), .Y(_19455_) );
	AOI21X1 AOI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_19454_), .B(_19432__bF_buf0), .C(_19455_), .Y(_17354__11_) );
	INVX1 INVX1_2827 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_12_), .Y(_19456_) );
	OAI21X1 OAI21X1_3906 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf60), .Y(_19457_) );
	AOI21X1 AOI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_19456_), .B(_19432__bF_buf6), .C(_19457_), .Y(_17354__12_) );
	INVX1 INVX1_2828 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_13_), .Y(_19458_) );
	OAI21X1 OAI21X1_3907 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf59), .Y(_19459_) );
	AOI21X1 AOI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_19458_), .B(_19432__bF_buf4), .C(_19459_), .Y(_17354__13_) );
	INVX1 INVX1_2829 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_14_), .Y(_19460_) );
	OAI21X1 OAI21X1_3908 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf58), .Y(_19461_) );
	AOI21X1 AOI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_19460_), .B(_19432__bF_buf2), .C(_19461_), .Y(_17354__14_) );
	INVX1 INVX1_2830 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_15_), .Y(_19462_) );
	OAI21X1 OAI21X1_3909 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf57), .Y(_19463_) );
	AOI21X1 AOI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_19462_), .B(_19432__bF_buf0), .C(_19463_), .Y(_17354__15_) );
	INVX1 INVX1_2831 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_16_), .Y(_19464_) );
	OAI21X1 OAI21X1_3910 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf56), .Y(_19465_) );
	AOI21X1 AOI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_19464_), .B(_19432__bF_buf6), .C(_19465_), .Y(_17354__16_) );
	INVX1 INVX1_2832 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_17_), .Y(_19466_) );
	OAI21X1 OAI21X1_3911 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf55), .Y(_19467_) );
	AOI21X1 AOI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_19466_), .B(_19432__bF_buf4), .C(_19467_), .Y(_17354__17_) );
	INVX1 INVX1_2833 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_18_), .Y(_19468_) );
	OAI21X1 OAI21X1_3912 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf54), .Y(_19469_) );
	AOI21X1 AOI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_19468_), .B(_19432__bF_buf2), .C(_19469_), .Y(_17354__18_) );
	INVX1 INVX1_2834 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_19_), .Y(_19470_) );
	OAI21X1 OAI21X1_3913 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf53), .Y(_19471_) );
	AOI21X1 AOI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_19470_), .B(_19432__bF_buf0), .C(_19471_), .Y(_17354__19_) );
	INVX1 INVX1_2835 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_20_), .Y(_19472_) );
	OAI21X1 OAI21X1_3914 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf52), .Y(_19473_) );
	AOI21X1 AOI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_19472_), .B(_19432__bF_buf6), .C(_19473_), .Y(_17354__20_) );
	INVX1 INVX1_2836 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_21_), .Y(_19474_) );
	OAI21X1 OAI21X1_3915 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf51), .Y(_19475_) );
	AOI21X1 AOI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_19474_), .B(_19432__bF_buf4), .C(_19475_), .Y(_17354__21_) );
	INVX1 INVX1_2837 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_22_), .Y(_19476_) );
	OAI21X1 OAI21X1_3916 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf50), .Y(_19477_) );
	AOI21X1 AOI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_19476_), .B(_19432__bF_buf2), .C(_19477_), .Y(_17354__22_) );
	INVX1 INVX1_2838 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_23_), .Y(_19478_) );
	OAI21X1 OAI21X1_3917 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf49), .Y(_19479_) );
	AOI21X1 AOI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_19478_), .B(_19432__bF_buf0), .C(_19479_), .Y(_17354__23_) );
	INVX1 INVX1_2839 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_24_), .Y(_19480_) );
	OAI21X1 OAI21X1_3918 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf48), .Y(_19481_) );
	AOI21X1 AOI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_19480_), .B(_19432__bF_buf6), .C(_19481_), .Y(_17354__24_) );
	INVX1 INVX1_2840 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_25_), .Y(_19482_) );
	OAI21X1 OAI21X1_3919 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf47), .Y(_19483_) );
	AOI21X1 AOI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_19482_), .B(_19432__bF_buf4), .C(_19483_), .Y(_17354__25_) );
	INVX1 INVX1_2841 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_26_), .Y(_19484_) );
	OAI21X1 OAI21X1_3920 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf46), .Y(_19485_) );
	AOI21X1 AOI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_19484_), .B(_19432__bF_buf2), .C(_19485_), .Y(_17354__26_) );
	INVX1 INVX1_2842 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_27_), .Y(_19486_) );
	OAI21X1 OAI21X1_3921 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf45), .Y(_19487_) );
	AOI21X1 AOI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_19486_), .B(_19432__bF_buf0), .C(_19487_), .Y(_17354__27_) );
	INVX1 INVX1_2843 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_28_), .Y(_19488_) );
	OAI21X1 OAI21X1_3922 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf2), .B(_19432__bF_buf7), .C(_19153__bF_buf44), .Y(_19489_) );
	AOI21X1 AOI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_19488_), .B(_19432__bF_buf6), .C(_19489_), .Y(_17354__28_) );
	INVX1 INVX1_2844 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_29_), .Y(_19490_) );
	OAI21X1 OAI21X1_3923 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf2), .B(_19432__bF_buf5), .C(_19153__bF_buf43), .Y(_19491_) );
	AOI21X1 AOI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_19490_), .B(_19432__bF_buf4), .C(_19491_), .Y(_17354__29_) );
	INVX1 INVX1_2845 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_30_), .Y(_19492_) );
	OAI21X1 OAI21X1_3924 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf2), .B(_19432__bF_buf3), .C(_19153__bF_buf42), .Y(_19493_) );
	AOI21X1 AOI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_19492_), .B(_19432__bF_buf2), .C(_19493_), .Y(_17354__30_) );
	INVX1 INVX1_2846 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_31_), .Y(_19494_) );
	OAI21X1 OAI21X1_3925 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf2), .B(_19432__bF_buf1), .C(_19153__bF_buf41), .Y(_19495_) );
	AOI21X1 AOI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_19494_), .B(_19432__bF_buf0), .C(_19495_), .Y(_17354__31_) );
	INVX1 INVX1_2847 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_3_), .Y(_19496_) );
	NAND2X1 NAND2X1_3550 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_2_), .B(_19496_), .Y(_19497_) );
	NOR2X1 NOR2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_19150_), .B(_19497_), .Y(_19498_) );
	NAND2X1 NAND2X1_3551 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19498_), .Y(_19499_) );
	OAI21X1 OAI21X1_3926 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf40), .Y(_19500_) );
	AOI21X1 AOI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_17448_), .B(_19499__bF_buf6), .C(_19500_), .Y(_17353__0_) );
	OAI21X1 OAI21X1_3927 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf39), .Y(_19501_) );
	AOI21X1 AOI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_17511_), .B(_19499__bF_buf4), .C(_19501_), .Y(_17353__1_) );
	OAI21X1 OAI21X1_3928 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf38), .Y(_19502_) );
	AOI21X1 AOI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_17565_), .B(_19499__bF_buf2), .C(_19502_), .Y(_17353__2_) );
	OAI21X1 OAI21X1_3929 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf37), .Y(_19503_) );
	AOI21X1 AOI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_17619_), .B(_19499__bF_buf0), .C(_19503_), .Y(_17353__3_) );
	OAI21X1 OAI21X1_3930 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf36), .Y(_19504_) );
	AOI21X1 AOI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_17673_), .B(_19499__bF_buf6), .C(_19504_), .Y(_17353__4_) );
	OAI21X1 OAI21X1_3931 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf35), .Y(_19505_) );
	AOI21X1 AOI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_17727_), .B(_19499__bF_buf4), .C(_19505_), .Y(_17353__5_) );
	OAI21X1 OAI21X1_3932 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf34), .Y(_19506_) );
	AOI21X1 AOI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_17781_), .B(_19499__bF_buf2), .C(_19506_), .Y(_17353__6_) );
	OAI21X1 OAI21X1_3933 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf33), .Y(_19507_) );
	AOI21X1 AOI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_17835_), .B(_19499__bF_buf0), .C(_19507_), .Y(_17353__7_) );
	OAI21X1 OAI21X1_3934 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf32), .Y(_19508_) );
	AOI21X1 AOI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_17889_), .B(_19499__bF_buf6), .C(_19508_), .Y(_17353__8_) );
	OAI21X1 OAI21X1_3935 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf31), .Y(_19509_) );
	AOI21X1 AOI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_17943_), .B(_19499__bF_buf4), .C(_19509_), .Y(_17353__9_) );
	OAI21X1 OAI21X1_3936 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf30), .Y(_19510_) );
	AOI21X1 AOI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_17997_), .B(_19499__bF_buf2), .C(_19510_), .Y(_17353__10_) );
	OAI21X1 OAI21X1_3937 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf29), .Y(_19511_) );
	AOI21X1 AOI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_18051_), .B(_19499__bF_buf0), .C(_19511_), .Y(_17353__11_) );
	OAI21X1 OAI21X1_3938 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf28), .Y(_19512_) );
	AOI21X1 AOI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_18105_), .B(_19499__bF_buf6), .C(_19512_), .Y(_17353__12_) );
	OAI21X1 OAI21X1_3939 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf27), .Y(_19513_) );
	AOI21X1 AOI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_18159_), .B(_19499__bF_buf4), .C(_19513_), .Y(_17353__13_) );
	OAI21X1 OAI21X1_3940 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf26), .Y(_19514_) );
	AOI21X1 AOI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_18213_), .B(_19499__bF_buf2), .C(_19514_), .Y(_17353__14_) );
	OAI21X1 OAI21X1_3941 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf25), .Y(_19515_) );
	AOI21X1 AOI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_18267_), .B(_19499__bF_buf0), .C(_19515_), .Y(_17353__15_) );
	OAI21X1 OAI21X1_3942 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf24), .Y(_19516_) );
	AOI21X1 AOI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_18321_), .B(_19499__bF_buf6), .C(_19516_), .Y(_17353__16_) );
	OAI21X1 OAI21X1_3943 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf23), .Y(_19517_) );
	AOI21X1 AOI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_18375_), .B(_19499__bF_buf4), .C(_19517_), .Y(_17353__17_) );
	OAI21X1 OAI21X1_3944 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf22), .Y(_19518_) );
	AOI21X1 AOI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_18429_), .B(_19499__bF_buf2), .C(_19518_), .Y(_17353__18_) );
	OAI21X1 OAI21X1_3945 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf21), .Y(_19519_) );
	AOI21X1 AOI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_18483_), .B(_19499__bF_buf0), .C(_19519_), .Y(_17353__19_) );
	OAI21X1 OAI21X1_3946 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf20), .Y(_19520_) );
	AOI21X1 AOI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_18537_), .B(_19499__bF_buf6), .C(_19520_), .Y(_17353__20_) );
	OAI21X1 OAI21X1_3947 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf19), .Y(_19521_) );
	AOI21X1 AOI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_18591_), .B(_19499__bF_buf4), .C(_19521_), .Y(_17353__21_) );
	OAI21X1 OAI21X1_3948 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf18), .Y(_19522_) );
	AOI21X1 AOI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_18645_), .B(_19499__bF_buf2), .C(_19522_), .Y(_17353__22_) );
	OAI21X1 OAI21X1_3949 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf17), .Y(_19523_) );
	AOI21X1 AOI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_18699_), .B(_19499__bF_buf0), .C(_19523_), .Y(_17353__23_) );
	OAI21X1 OAI21X1_3950 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf16), .Y(_19524_) );
	AOI21X1 AOI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_18753_), .B(_19499__bF_buf6), .C(_19524_), .Y(_17353__24_) );
	OAI21X1 OAI21X1_3951 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf15), .Y(_19525_) );
	AOI21X1 AOI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_18807_), .B(_19499__bF_buf4), .C(_19525_), .Y(_17353__25_) );
	OAI21X1 OAI21X1_3952 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf14), .Y(_19526_) );
	AOI21X1 AOI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_18861_), .B(_19499__bF_buf2), .C(_19526_), .Y(_17353__26_) );
	OAI21X1 OAI21X1_3953 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf13), .Y(_19527_) );
	AOI21X1 AOI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_18915_), .B(_19499__bF_buf0), .C(_19527_), .Y(_17353__27_) );
	OAI21X1 OAI21X1_3954 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf1), .B(_19499__bF_buf7), .C(_19153__bF_buf12), .Y(_19528_) );
	AOI21X1 AOI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_18969_), .B(_19499__bF_buf6), .C(_19528_), .Y(_17353__28_) );
	OAI21X1 OAI21X1_3955 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf1), .B(_19499__bF_buf5), .C(_19153__bF_buf11), .Y(_19529_) );
	AOI21X1 AOI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_19023_), .B(_19499__bF_buf4), .C(_19529_), .Y(_17353__29_) );
	OAI21X1 OAI21X1_3956 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf1), .B(_19499__bF_buf3), .C(_19153__bF_buf10), .Y(_19530_) );
	AOI21X1 AOI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_19077_), .B(_19499__bF_buf2), .C(_19530_), .Y(_17353__30_) );
	OAI21X1 OAI21X1_3957 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf1), .B(_19499__bF_buf1), .C(_19153__bF_buf9), .Y(_19531_) );
	AOI21X1 AOI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_19131_), .B(_19499__bF_buf0), .C(_19531_), .Y(_17353__31_) );
	NOR2X1 NOR2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_19218_), .B(_19497_), .Y(_19532_) );
	NAND2X1 NAND2X1_3552 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19532_), .Y(_19533_) );
	OAI21X1 OAI21X1_3958 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf8), .Y(_19534_) );
	AOI21X1 AOI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_17447_), .B(_19533__bF_buf6), .C(_19534_), .Y(_17352__0_) );
	OAI21X1 OAI21X1_3959 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf7), .Y(_19535_) );
	AOI21X1 AOI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_17510_), .B(_19533__bF_buf4), .C(_19535_), .Y(_17352__1_) );
	OAI21X1 OAI21X1_3960 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf6), .Y(_19536_) );
	AOI21X1 AOI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_17564_), .B(_19533__bF_buf2), .C(_19536_), .Y(_17352__2_) );
	OAI21X1 OAI21X1_3961 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf5), .Y(_19537_) );
	AOI21X1 AOI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_17618_), .B(_19533__bF_buf0), .C(_19537_), .Y(_17352__3_) );
	OAI21X1 OAI21X1_3962 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf4), .Y(_19538_) );
	AOI21X1 AOI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_17672_), .B(_19533__bF_buf6), .C(_19538_), .Y(_17352__4_) );
	OAI21X1 OAI21X1_3963 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf3), .Y(_19539_) );
	AOI21X1 AOI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_17726_), .B(_19533__bF_buf4), .C(_19539_), .Y(_17352__5_) );
	OAI21X1 OAI21X1_3964 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf2), .Y(_19540_) );
	AOI21X1 AOI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_17780_), .B(_19533__bF_buf2), .C(_19540_), .Y(_17352__6_) );
	OAI21X1 OAI21X1_3965 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf1), .Y(_19541_) );
	AOI21X1 AOI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_17834_), .B(_19533__bF_buf0), .C(_19541_), .Y(_17352__7_) );
	OAI21X1 OAI21X1_3966 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf0), .Y(_19542_) );
	AOI21X1 AOI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_17888_), .B(_19533__bF_buf6), .C(_19542_), .Y(_17352__8_) );
	OAI21X1 OAI21X1_3967 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf98), .Y(_19543_) );
	AOI21X1 AOI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_17942_), .B(_19533__bF_buf4), .C(_19543_), .Y(_17352__9_) );
	OAI21X1 OAI21X1_3968 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf97), .Y(_19544_) );
	AOI21X1 AOI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_17996_), .B(_19533__bF_buf2), .C(_19544_), .Y(_17352__10_) );
	OAI21X1 OAI21X1_3969 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf96), .Y(_19545_) );
	AOI21X1 AOI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_18050_), .B(_19533__bF_buf0), .C(_19545_), .Y(_17352__11_) );
	OAI21X1 OAI21X1_3970 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf95), .Y(_19546_) );
	AOI21X1 AOI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_18104_), .B(_19533__bF_buf6), .C(_19546_), .Y(_17352__12_) );
	OAI21X1 OAI21X1_3971 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf94), .Y(_19547_) );
	AOI21X1 AOI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_18158_), .B(_19533__bF_buf4), .C(_19547_), .Y(_17352__13_) );
	OAI21X1 OAI21X1_3972 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf93), .Y(_19548_) );
	AOI21X1 AOI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_18212_), .B(_19533__bF_buf2), .C(_19548_), .Y(_17352__14_) );
	OAI21X1 OAI21X1_3973 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf92), .Y(_19549_) );
	AOI21X1 AOI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_18266_), .B(_19533__bF_buf0), .C(_19549_), .Y(_17352__15_) );
	OAI21X1 OAI21X1_3974 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf91), .Y(_19550_) );
	AOI21X1 AOI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_18320_), .B(_19533__bF_buf6), .C(_19550_), .Y(_17352__16_) );
	OAI21X1 OAI21X1_3975 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf90), .Y(_19551_) );
	AOI21X1 AOI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_18374_), .B(_19533__bF_buf4), .C(_19551_), .Y(_17352__17_) );
	OAI21X1 OAI21X1_3976 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf89), .Y(_19552_) );
	AOI21X1 AOI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_18428_), .B(_19533__bF_buf2), .C(_19552_), .Y(_17352__18_) );
	OAI21X1 OAI21X1_3977 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf88), .Y(_19553_) );
	AOI21X1 AOI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_18482_), .B(_19533__bF_buf0), .C(_19553_), .Y(_17352__19_) );
	OAI21X1 OAI21X1_3978 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf87), .Y(_19554_) );
	AOI21X1 AOI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_18536_), .B(_19533__bF_buf6), .C(_19554_), .Y(_17352__20_) );
	OAI21X1 OAI21X1_3979 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf86), .Y(_19555_) );
	AOI21X1 AOI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_18590_), .B(_19533__bF_buf4), .C(_19555_), .Y(_17352__21_) );
	OAI21X1 OAI21X1_3980 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf85), .Y(_19556_) );
	AOI21X1 AOI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_18644_), .B(_19533__bF_buf2), .C(_19556_), .Y(_17352__22_) );
	OAI21X1 OAI21X1_3981 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf84), .Y(_19557_) );
	AOI21X1 AOI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_18698_), .B(_19533__bF_buf0), .C(_19557_), .Y(_17352__23_) );
	OAI21X1 OAI21X1_3982 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf83), .Y(_19558_) );
	AOI21X1 AOI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_18752_), .B(_19533__bF_buf6), .C(_19558_), .Y(_17352__24_) );
	OAI21X1 OAI21X1_3983 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf82), .Y(_19559_) );
	AOI21X1 AOI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_18806_), .B(_19533__bF_buf4), .C(_19559_), .Y(_17352__25_) );
	OAI21X1 OAI21X1_3984 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf81), .Y(_19560_) );
	AOI21X1 AOI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_18860_), .B(_19533__bF_buf2), .C(_19560_), .Y(_17352__26_) );
	OAI21X1 OAI21X1_3985 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf80), .Y(_19561_) );
	AOI21X1 AOI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_18914_), .B(_19533__bF_buf0), .C(_19561_), .Y(_17352__27_) );
	OAI21X1 OAI21X1_3986 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf0), .B(_19533__bF_buf7), .C(_19153__bF_buf79), .Y(_19562_) );
	AOI21X1 AOI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_18968_), .B(_19533__bF_buf6), .C(_19562_), .Y(_17352__28_) );
	OAI21X1 OAI21X1_3987 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf0), .B(_19533__bF_buf5), .C(_19153__bF_buf78), .Y(_19563_) );
	AOI21X1 AOI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_19022_), .B(_19533__bF_buf4), .C(_19563_), .Y(_17352__29_) );
	OAI21X1 OAI21X1_3988 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf0), .B(_19533__bF_buf3), .C(_19153__bF_buf77), .Y(_19564_) );
	AOI21X1 AOI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_19076_), .B(_19533__bF_buf2), .C(_19564_), .Y(_17352__30_) );
	OAI21X1 OAI21X1_3989 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf0), .B(_19533__bF_buf1), .C(_19153__bF_buf76), .Y(_19565_) );
	AOI21X1 AOI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_19130_), .B(_19533__bF_buf0), .C(_19565_), .Y(_17352__31_) );
	NOR2X1 NOR2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_19254_), .B(_19497_), .Y(_19566_) );
	NAND2X1 NAND2X1_3553 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19566_), .Y(_19567_) );
	OAI21X1 OAI21X1_3990 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf75), .Y(_19568_) );
	AOI21X1 AOI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_17410_), .B(_19567__bF_buf6), .C(_19568_), .Y(_17351__0_) );
	OAI21X1 OAI21X1_3991 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf74), .Y(_19569_) );
	AOI21X1 AOI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_17490_), .B(_19567__bF_buf4), .C(_19569_), .Y(_17351__1_) );
	OAI21X1 OAI21X1_3992 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf73), .Y(_19570_) );
	AOI21X1 AOI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_17544_), .B(_19567__bF_buf2), .C(_19570_), .Y(_17351__2_) );
	OAI21X1 OAI21X1_3993 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf72), .Y(_19571_) );
	AOI21X1 AOI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_17598_), .B(_19567__bF_buf0), .C(_19571_), .Y(_17351__3_) );
	OAI21X1 OAI21X1_3994 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf71), .Y(_19572_) );
	AOI21X1 AOI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_17652_), .B(_19567__bF_buf6), .C(_19572_), .Y(_17351__4_) );
	OAI21X1 OAI21X1_3995 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf70), .Y(_19573_) );
	AOI21X1 AOI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_17706_), .B(_19567__bF_buf4), .C(_19573_), .Y(_17351__5_) );
	OAI21X1 OAI21X1_3996 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf69), .Y(_19574_) );
	AOI21X1 AOI21X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_17760_), .B(_19567__bF_buf2), .C(_19574_), .Y(_17351__6_) );
	OAI21X1 OAI21X1_3997 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf68), .Y(_19575_) );
	AOI21X1 AOI21X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_17814_), .B(_19567__bF_buf0), .C(_19575_), .Y(_17351__7_) );
	OAI21X1 OAI21X1_3998 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf67), .Y(_19576_) );
	AOI21X1 AOI21X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_17868_), .B(_19567__bF_buf6), .C(_19576_), .Y(_17351__8_) );
	OAI21X1 OAI21X1_3999 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf66), .Y(_19577_) );
	AOI21X1 AOI21X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_17922_), .B(_19567__bF_buf4), .C(_19577_), .Y(_17351__9_) );
	OAI21X1 OAI21X1_4000 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf65), .Y(_19578_) );
	AOI21X1 AOI21X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_17976_), .B(_19567__bF_buf2), .C(_19578_), .Y(_17351__10_) );
	OAI21X1 OAI21X1_4001 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf64), .Y(_19579_) );
	AOI21X1 AOI21X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_18030_), .B(_19567__bF_buf0), .C(_19579_), .Y(_17351__11_) );
	OAI21X1 OAI21X1_4002 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf63), .Y(_19580_) );
	AOI21X1 AOI21X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_18084_), .B(_19567__bF_buf6), .C(_19580_), .Y(_17351__12_) );
	OAI21X1 OAI21X1_4003 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf62), .Y(_19581_) );
	AOI21X1 AOI21X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_18138_), .B(_19567__bF_buf4), .C(_19581_), .Y(_17351__13_) );
	OAI21X1 OAI21X1_4004 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf61), .Y(_19582_) );
	AOI21X1 AOI21X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_18192_), .B(_19567__bF_buf2), .C(_19582_), .Y(_17351__14_) );
	OAI21X1 OAI21X1_4005 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf60), .Y(_19583_) );
	AOI21X1 AOI21X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_18246_), .B(_19567__bF_buf0), .C(_19583_), .Y(_17351__15_) );
	OAI21X1 OAI21X1_4006 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf59), .Y(_19584_) );
	AOI21X1 AOI21X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_18300_), .B(_19567__bF_buf6), .C(_19584_), .Y(_17351__16_) );
	OAI21X1 OAI21X1_4007 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf58), .Y(_19585_) );
	AOI21X1 AOI21X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_18354_), .B(_19567__bF_buf4), .C(_19585_), .Y(_17351__17_) );
	OAI21X1 OAI21X1_4008 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf57), .Y(_19586_) );
	AOI21X1 AOI21X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_18408_), .B(_19567__bF_buf2), .C(_19586_), .Y(_17351__18_) );
	OAI21X1 OAI21X1_4009 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf56), .Y(_19587_) );
	AOI21X1 AOI21X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_18462_), .B(_19567__bF_buf0), .C(_19587_), .Y(_17351__19_) );
	OAI21X1 OAI21X1_4010 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf55), .Y(_19588_) );
	AOI21X1 AOI21X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_18516_), .B(_19567__bF_buf6), .C(_19588_), .Y(_17351__20_) );
	OAI21X1 OAI21X1_4011 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf54), .Y(_19589_) );
	AOI21X1 AOI21X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_18570_), .B(_19567__bF_buf4), .C(_19589_), .Y(_17351__21_) );
	OAI21X1 OAI21X1_4012 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf53), .Y(_19590_) );
	AOI21X1 AOI21X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_18624_), .B(_19567__bF_buf2), .C(_19590_), .Y(_17351__22_) );
	OAI21X1 OAI21X1_4013 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf52), .Y(_19591_) );
	AOI21X1 AOI21X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_18678_), .B(_19567__bF_buf0), .C(_19591_), .Y(_17351__23_) );
	OAI21X1 OAI21X1_4014 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf51), .Y(_19592_) );
	AOI21X1 AOI21X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_18732_), .B(_19567__bF_buf6), .C(_19592_), .Y(_17351__24_) );
	OAI21X1 OAI21X1_4015 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf50), .Y(_19593_) );
	AOI21X1 AOI21X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_18786_), .B(_19567__bF_buf4), .C(_19593_), .Y(_17351__25_) );
	OAI21X1 OAI21X1_4016 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf49), .Y(_19594_) );
	AOI21X1 AOI21X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_18840_), .B(_19567__bF_buf2), .C(_19594_), .Y(_17351__26_) );
	OAI21X1 OAI21X1_4017 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf48), .Y(_19595_) );
	AOI21X1 AOI21X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_18894_), .B(_19567__bF_buf0), .C(_19595_), .Y(_17351__27_) );
	OAI21X1 OAI21X1_4018 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_19567__bF_buf7), .C(_19153__bF_buf47), .Y(_19596_) );
	AOI21X1 AOI21X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_18948_), .B(_19567__bF_buf6), .C(_19596_), .Y(_17351__28_) );
	OAI21X1 OAI21X1_4019 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_19567__bF_buf5), .C(_19153__bF_buf46), .Y(_19597_) );
	AOI21X1 AOI21X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_19002_), .B(_19567__bF_buf4), .C(_19597_), .Y(_17351__29_) );
	OAI21X1 OAI21X1_4020 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_19567__bF_buf3), .C(_19153__bF_buf45), .Y(_19598_) );
	AOI21X1 AOI21X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_19056_), .B(_19567__bF_buf2), .C(_19598_), .Y(_17351__30_) );
	OAI21X1 OAI21X1_4021 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_19567__bF_buf1), .C(_19153__bF_buf44), .Y(_19599_) );
	AOI21X1 AOI21X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_19110_), .B(_19567__bF_buf0), .C(_19599_), .Y(_17351__31_) );
	INVX1 INVX1_2848 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_0_), .Y(_19600_) );
	INVX1 INVX1_2849 ( .gnd(gnd), .vdd(vdd), .A(_19497_), .Y(_19601_) );
	NAND2X1 NAND2X1_3554 ( .gnd(gnd), .vdd(vdd), .A(_19601_), .B(_19430_), .Y(_19602_) );
	OAI21X1 OAI21X1_4022 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf43), .Y(_19603_) );
	AOI21X1 AOI21X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_19600_), .B(_19602__bF_buf6), .C(_19603_), .Y(_17350__0_) );
	INVX1 INVX1_2850 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_1_), .Y(_19604_) );
	OAI21X1 OAI21X1_4023 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf42), .Y(_19605_) );
	AOI21X1 AOI21X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_19604_), .B(_19602__bF_buf4), .C(_19605_), .Y(_17350__1_) );
	INVX1 INVX1_2851 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_2_), .Y(_19606_) );
	OAI21X1 OAI21X1_4024 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf41), .Y(_19607_) );
	AOI21X1 AOI21X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_19606_), .B(_19602__bF_buf2), .C(_19607_), .Y(_17350__2_) );
	INVX1 INVX1_2852 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_3_), .Y(_19608_) );
	OAI21X1 OAI21X1_4025 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf40), .Y(_19609_) );
	AOI21X1 AOI21X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_19608_), .B(_19602__bF_buf0), .C(_19609_), .Y(_17350__3_) );
	INVX1 INVX1_2853 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_4_), .Y(_19610_) );
	OAI21X1 OAI21X1_4026 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf39), .Y(_19611_) );
	AOI21X1 AOI21X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_19610_), .B(_19602__bF_buf6), .C(_19611_), .Y(_17350__4_) );
	INVX1 INVX1_2854 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_5_), .Y(_19612_) );
	OAI21X1 OAI21X1_4027 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf38), .Y(_19613_) );
	AOI21X1 AOI21X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_19612_), .B(_19602__bF_buf4), .C(_19613_), .Y(_17350__5_) );
	INVX1 INVX1_2855 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_6_), .Y(_19614_) );
	OAI21X1 OAI21X1_4028 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf37), .Y(_19615_) );
	AOI21X1 AOI21X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_19614_), .B(_19602__bF_buf2), .C(_19615_), .Y(_17350__6_) );
	INVX1 INVX1_2856 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_7_), .Y(_19616_) );
	OAI21X1 OAI21X1_4029 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf36), .Y(_19617_) );
	AOI21X1 AOI21X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_19616_), .B(_19602__bF_buf0), .C(_19617_), .Y(_17350__7_) );
	INVX1 INVX1_2857 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_8_), .Y(_19618_) );
	OAI21X1 OAI21X1_4030 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf35), .Y(_19619_) );
	AOI21X1 AOI21X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_19618_), .B(_19602__bF_buf6), .C(_19619_), .Y(_17350__8_) );
	INVX1 INVX1_2858 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_9_), .Y(_19620_) );
	OAI21X1 OAI21X1_4031 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf34), .Y(_19621_) );
	AOI21X1 AOI21X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_19620_), .B(_19602__bF_buf4), .C(_19621_), .Y(_17350__9_) );
	INVX1 INVX1_2859 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_10_), .Y(_19622_) );
	OAI21X1 OAI21X1_4032 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf33), .Y(_19623_) );
	AOI21X1 AOI21X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_19622_), .B(_19602__bF_buf2), .C(_19623_), .Y(_17350__10_) );
	INVX1 INVX1_2860 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_11_), .Y(_19624_) );
	OAI21X1 OAI21X1_4033 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf32), .Y(_19625_) );
	AOI21X1 AOI21X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_19624_), .B(_19602__bF_buf0), .C(_19625_), .Y(_17350__11_) );
	INVX1 INVX1_2861 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_12_), .Y(_19626_) );
	OAI21X1 OAI21X1_4034 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf31), .Y(_19627_) );
	AOI21X1 AOI21X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_19626_), .B(_19602__bF_buf6), .C(_19627_), .Y(_17350__12_) );
	INVX1 INVX1_2862 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_13_), .Y(_19628_) );
	OAI21X1 OAI21X1_4035 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf30), .Y(_19629_) );
	AOI21X1 AOI21X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_19628_), .B(_19602__bF_buf4), .C(_19629_), .Y(_17350__13_) );
	INVX1 INVX1_2863 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_14_), .Y(_19630_) );
	OAI21X1 OAI21X1_4036 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf29), .Y(_19631_) );
	AOI21X1 AOI21X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_19630_), .B(_19602__bF_buf2), .C(_19631_), .Y(_17350__14_) );
	INVX1 INVX1_2864 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_15_), .Y(_19632_) );
	OAI21X1 OAI21X1_4037 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf28), .Y(_19633_) );
	AOI21X1 AOI21X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_19632_), .B(_19602__bF_buf0), .C(_19633_), .Y(_17350__15_) );
	INVX1 INVX1_2865 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_16_), .Y(_19634_) );
	OAI21X1 OAI21X1_4038 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf27), .Y(_19635_) );
	AOI21X1 AOI21X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_19634_), .B(_19602__bF_buf6), .C(_19635_), .Y(_17350__16_) );
	INVX1 INVX1_2866 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_17_), .Y(_19636_) );
	OAI21X1 OAI21X1_4039 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf26), .Y(_19637_) );
	AOI21X1 AOI21X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_19636_), .B(_19602__bF_buf4), .C(_19637_), .Y(_17350__17_) );
	INVX1 INVX1_2867 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_18_), .Y(_19638_) );
	OAI21X1 OAI21X1_4040 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf25), .Y(_19639_) );
	AOI21X1 AOI21X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_19638_), .B(_19602__bF_buf2), .C(_19639_), .Y(_17350__18_) );
	INVX1 INVX1_2868 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_19_), .Y(_19640_) );
	OAI21X1 OAI21X1_4041 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf24), .Y(_19641_) );
	AOI21X1 AOI21X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_19640_), .B(_19602__bF_buf0), .C(_19641_), .Y(_17350__19_) );
	INVX1 INVX1_2869 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_20_), .Y(_19642_) );
	OAI21X1 OAI21X1_4042 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf23), .Y(_19643_) );
	AOI21X1 AOI21X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_19642_), .B(_19602__bF_buf6), .C(_19643_), .Y(_17350__20_) );
	INVX1 INVX1_2870 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_21_), .Y(_19644_) );
	OAI21X1 OAI21X1_4043 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf22), .Y(_19645_) );
	AOI21X1 AOI21X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_19644_), .B(_19602__bF_buf4), .C(_19645_), .Y(_17350__21_) );
	INVX1 INVX1_2871 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_22_), .Y(_19646_) );
	OAI21X1 OAI21X1_4044 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf21), .Y(_19647_) );
	AOI21X1 AOI21X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_19646_), .B(_19602__bF_buf2), .C(_19647_), .Y(_17350__22_) );
	INVX1 INVX1_2872 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_23_), .Y(_19648_) );
	OAI21X1 OAI21X1_4045 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf20), .Y(_19649_) );
	AOI21X1 AOI21X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_19648_), .B(_19602__bF_buf0), .C(_19649_), .Y(_17350__23_) );
	INVX1 INVX1_2873 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_24_), .Y(_19650_) );
	OAI21X1 OAI21X1_4046 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf19), .Y(_19651_) );
	AOI21X1 AOI21X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_19650_), .B(_19602__bF_buf6), .C(_19651_), .Y(_17350__24_) );
	INVX1 INVX1_2874 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_25_), .Y(_19652_) );
	OAI21X1 OAI21X1_4047 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf18), .Y(_19653_) );
	AOI21X1 AOI21X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_19652_), .B(_19602__bF_buf4), .C(_19653_), .Y(_17350__25_) );
	INVX1 INVX1_2875 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_26_), .Y(_19654_) );
	OAI21X1 OAI21X1_4048 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf17), .Y(_19655_) );
	AOI21X1 AOI21X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_19654_), .B(_19602__bF_buf2), .C(_19655_), .Y(_17350__26_) );
	INVX1 INVX1_2876 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_27_), .Y(_19656_) );
	OAI21X1 OAI21X1_4049 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf16), .Y(_19657_) );
	AOI21X1 AOI21X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_19656_), .B(_19602__bF_buf0), .C(_19657_), .Y(_17350__27_) );
	INVX1 INVX1_2877 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_28_), .Y(_19658_) );
	OAI21X1 OAI21X1_4050 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf3), .B(_19602__bF_buf7), .C(_19153__bF_buf15), .Y(_19659_) );
	AOI21X1 AOI21X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_19658_), .B(_19602__bF_buf6), .C(_19659_), .Y(_17350__28_) );
	INVX1 INVX1_2878 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_29_), .Y(_19660_) );
	OAI21X1 OAI21X1_4051 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf3), .B(_19602__bF_buf5), .C(_19153__bF_buf14), .Y(_19661_) );
	AOI21X1 AOI21X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_19660_), .B(_19602__bF_buf4), .C(_19661_), .Y(_17350__29_) );
	INVX1 INVX1_2879 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_30_), .Y(_19662_) );
	OAI21X1 OAI21X1_4052 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf3), .B(_19602__bF_buf3), .C(_19153__bF_buf13), .Y(_19663_) );
	AOI21X1 AOI21X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_19662_), .B(_19602__bF_buf2), .C(_19663_), .Y(_17350__30_) );
	INVX1 INVX1_2880 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_31_), .Y(_19664_) );
	OAI21X1 OAI21X1_4053 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf3), .B(_19602__bF_buf1), .C(_19153__bF_buf12), .Y(_19665_) );
	AOI21X1 AOI21X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_19664_), .B(_19602__bF_buf0), .C(_19665_), .Y(_17350__31_) );
	NAND2X1 NAND2X1_3555 ( .gnd(gnd), .vdd(vdd), .A(_19496_), .B(_19325_), .Y(_19666_) );
	NOR2X1 NOR2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_19150_), .B(_19666_), .Y(_19667_) );
	NAND2X1 NAND2X1_3556 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19667_), .Y(_19668_) );
	OAI21X1 OAI21X1_4054 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf11), .Y(_19669_) );
	AOI21X1 AOI21X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_17406_), .B(_19668__bF_buf6), .C(_19669_), .Y(_17348__0_) );
	OAI21X1 OAI21X1_4055 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf10), .Y(_19670_) );
	AOI21X1 AOI21X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_17488_), .B(_19668__bF_buf4), .C(_19670_), .Y(_17348__1_) );
	OAI21X1 OAI21X1_4056 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf9), .Y(_19671_) );
	AOI21X1 AOI21X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_17542_), .B(_19668__bF_buf2), .C(_19671_), .Y(_17348__2_) );
	OAI21X1 OAI21X1_4057 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf8), .Y(_19672_) );
	AOI21X1 AOI21X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_17596_), .B(_19668__bF_buf0), .C(_19672_), .Y(_17348__3_) );
	OAI21X1 OAI21X1_4058 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf7), .Y(_19673_) );
	AOI21X1 AOI21X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_17650_), .B(_19668__bF_buf6), .C(_19673_), .Y(_17348__4_) );
	OAI21X1 OAI21X1_4059 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf6), .Y(_19674_) );
	AOI21X1 AOI21X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_17704_), .B(_19668__bF_buf4), .C(_19674_), .Y(_17348__5_) );
	OAI21X1 OAI21X1_4060 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf5), .Y(_19675_) );
	AOI21X1 AOI21X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_17758_), .B(_19668__bF_buf2), .C(_19675_), .Y(_17348__6_) );
	OAI21X1 OAI21X1_4061 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf4), .Y(_19676_) );
	AOI21X1 AOI21X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_17812_), .B(_19668__bF_buf0), .C(_19676_), .Y(_17348__7_) );
	OAI21X1 OAI21X1_4062 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf3), .Y(_19677_) );
	AOI21X1 AOI21X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_17866_), .B(_19668__bF_buf6), .C(_19677_), .Y(_17348__8_) );
	OAI21X1 OAI21X1_4063 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf2), .Y(_19678_) );
	AOI21X1 AOI21X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_17920_), .B(_19668__bF_buf4), .C(_19678_), .Y(_17348__9_) );
	OAI21X1 OAI21X1_4064 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf1), .Y(_19679_) );
	AOI21X1 AOI21X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_17974_), .B(_19668__bF_buf2), .C(_19679_), .Y(_17348__10_) );
	OAI21X1 OAI21X1_4065 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf0), .Y(_19680_) );
	AOI21X1 AOI21X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_18028_), .B(_19668__bF_buf0), .C(_19680_), .Y(_17348__11_) );
	OAI21X1 OAI21X1_4066 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf98), .Y(_19681_) );
	AOI21X1 AOI21X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_18082_), .B(_19668__bF_buf6), .C(_19681_), .Y(_17348__12_) );
	OAI21X1 OAI21X1_4067 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf97), .Y(_19682_) );
	AOI21X1 AOI21X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_18136_), .B(_19668__bF_buf4), .C(_19682_), .Y(_17348__13_) );
	OAI21X1 OAI21X1_4068 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf96), .Y(_19683_) );
	AOI21X1 AOI21X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_18190_), .B(_19668__bF_buf2), .C(_19683_), .Y(_17348__14_) );
	OAI21X1 OAI21X1_4069 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf95), .Y(_19684_) );
	AOI21X1 AOI21X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_18244_), .B(_19668__bF_buf0), .C(_19684_), .Y(_17348__15_) );
	OAI21X1 OAI21X1_4070 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf94), .Y(_19685_) );
	AOI21X1 AOI21X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_18298_), .B(_19668__bF_buf6), .C(_19685_), .Y(_17348__16_) );
	OAI21X1 OAI21X1_4071 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf93), .Y(_19686_) );
	AOI21X1 AOI21X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_18352_), .B(_19668__bF_buf4), .C(_19686_), .Y(_17348__17_) );
	OAI21X1 OAI21X1_4072 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf92), .Y(_19687_) );
	AOI21X1 AOI21X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_18406_), .B(_19668__bF_buf2), .C(_19687_), .Y(_17348__18_) );
	OAI21X1 OAI21X1_4073 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf91), .Y(_19688_) );
	AOI21X1 AOI21X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_18460_), .B(_19668__bF_buf0), .C(_19688_), .Y(_17348__19_) );
	OAI21X1 OAI21X1_4074 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf90), .Y(_19689_) );
	AOI21X1 AOI21X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_18514_), .B(_19668__bF_buf6), .C(_19689_), .Y(_17348__20_) );
	OAI21X1 OAI21X1_4075 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf89), .Y(_19690_) );
	AOI21X1 AOI21X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_18568_), .B(_19668__bF_buf4), .C(_19690_), .Y(_17348__21_) );
	OAI21X1 OAI21X1_4076 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf88), .Y(_19691_) );
	AOI21X1 AOI21X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_18622_), .B(_19668__bF_buf2), .C(_19691_), .Y(_17348__22_) );
	OAI21X1 OAI21X1_4077 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf87), .Y(_19692_) );
	AOI21X1 AOI21X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_18676_), .B(_19668__bF_buf0), .C(_19692_), .Y(_17348__23_) );
	OAI21X1 OAI21X1_4078 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf86), .Y(_19693_) );
	AOI21X1 AOI21X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_18730_), .B(_19668__bF_buf6), .C(_19693_), .Y(_17348__24_) );
	OAI21X1 OAI21X1_4079 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf85), .Y(_19694_) );
	AOI21X1 AOI21X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_18784_), .B(_19668__bF_buf4), .C(_19694_), .Y(_17348__25_) );
	OAI21X1 OAI21X1_4080 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf84), .Y(_19695_) );
	AOI21X1 AOI21X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_18838_), .B(_19668__bF_buf2), .C(_19695_), .Y(_17348__26_) );
	OAI21X1 OAI21X1_4081 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf83), .Y(_19696_) );
	AOI21X1 AOI21X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_18892_), .B(_19668__bF_buf0), .C(_19696_), .Y(_17348__27_) );
	OAI21X1 OAI21X1_4082 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf2), .B(_19668__bF_buf7), .C(_19153__bF_buf82), .Y(_19697_) );
	AOI21X1 AOI21X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_18946_), .B(_19668__bF_buf6), .C(_19697_), .Y(_17348__28_) );
	OAI21X1 OAI21X1_4083 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf2), .B(_19668__bF_buf5), .C(_19153__bF_buf81), .Y(_19698_) );
	AOI21X1 AOI21X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_19000_), .B(_19668__bF_buf4), .C(_19698_), .Y(_17348__29_) );
	OAI21X1 OAI21X1_4084 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf2), .B(_19668__bF_buf3), .C(_19153__bF_buf80), .Y(_19699_) );
	AOI21X1 AOI21X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_19054_), .B(_19668__bF_buf2), .C(_19699_), .Y(_17348__30_) );
	OAI21X1 OAI21X1_4085 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf2), .B(_19668__bF_buf1), .C(_19153__bF_buf79), .Y(_19700_) );
	AOI21X1 AOI21X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_19108_), .B(_19668__bF_buf0), .C(_19700_), .Y(_17348__31_) );
	NOR2X1 NOR2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_19218_), .B(_19666_), .Y(_19701_) );
	NAND2X1 NAND2X1_3557 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19701_), .Y(_19702_) );
	OAI21X1 OAI21X1_4086 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf78), .Y(_19703_) );
	AOI21X1 AOI21X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_17405_), .B(_19702__bF_buf6), .C(_19703_), .Y(_17347__0_) );
	OAI21X1 OAI21X1_4087 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf77), .Y(_19704_) );
	AOI21X1 AOI21X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_17487_), .B(_19702__bF_buf4), .C(_19704_), .Y(_17347__1_) );
	OAI21X1 OAI21X1_4088 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf76), .Y(_19705_) );
	AOI21X1 AOI21X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_17541_), .B(_19702__bF_buf2), .C(_19705_), .Y(_17347__2_) );
	OAI21X1 OAI21X1_4089 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf75), .Y(_19706_) );
	AOI21X1 AOI21X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_17595_), .B(_19702__bF_buf0), .C(_19706_), .Y(_17347__3_) );
	OAI21X1 OAI21X1_4090 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf74), .Y(_19707_) );
	AOI21X1 AOI21X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_17649_), .B(_19702__bF_buf6), .C(_19707_), .Y(_17347__4_) );
	OAI21X1 OAI21X1_4091 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf73), .Y(_19708_) );
	AOI21X1 AOI21X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_17703_), .B(_19702__bF_buf4), .C(_19708_), .Y(_17347__5_) );
	OAI21X1 OAI21X1_4092 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf72), .Y(_19709_) );
	AOI21X1 AOI21X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_17757_), .B(_19702__bF_buf2), .C(_19709_), .Y(_17347__6_) );
	OAI21X1 OAI21X1_4093 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf71), .Y(_19710_) );
	AOI21X1 AOI21X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_17811_), .B(_19702__bF_buf0), .C(_19710_), .Y(_17347__7_) );
	OAI21X1 OAI21X1_4094 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf70), .Y(_19711_) );
	AOI21X1 AOI21X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_17865_), .B(_19702__bF_buf6), .C(_19711_), .Y(_17347__8_) );
	OAI21X1 OAI21X1_4095 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf69), .Y(_19712_) );
	AOI21X1 AOI21X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_17919_), .B(_19702__bF_buf4), .C(_19712_), .Y(_17347__9_) );
	OAI21X1 OAI21X1_4096 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf68), .Y(_19713_) );
	AOI21X1 AOI21X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_17973_), .B(_19702__bF_buf2), .C(_19713_), .Y(_17347__10_) );
	OAI21X1 OAI21X1_4097 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf67), .Y(_19714_) );
	AOI21X1 AOI21X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_18027_), .B(_19702__bF_buf0), .C(_19714_), .Y(_17347__11_) );
	OAI21X1 OAI21X1_4098 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf66), .Y(_19715_) );
	AOI21X1 AOI21X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_18081_), .B(_19702__bF_buf6), .C(_19715_), .Y(_17347__12_) );
	OAI21X1 OAI21X1_4099 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf65), .Y(_19716_) );
	AOI21X1 AOI21X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_18135_), .B(_19702__bF_buf4), .C(_19716_), .Y(_17347__13_) );
	OAI21X1 OAI21X1_4100 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf64), .Y(_19717_) );
	AOI21X1 AOI21X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_18189_), .B(_19702__bF_buf2), .C(_19717_), .Y(_17347__14_) );
	OAI21X1 OAI21X1_4101 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf63), .Y(_19718_) );
	AOI21X1 AOI21X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_18243_), .B(_19702__bF_buf0), .C(_19718_), .Y(_17347__15_) );
	OAI21X1 OAI21X1_4102 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf62), .Y(_19719_) );
	AOI21X1 AOI21X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_18297_), .B(_19702__bF_buf6), .C(_19719_), .Y(_17347__16_) );
	OAI21X1 OAI21X1_4103 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf61), .Y(_19720_) );
	AOI21X1 AOI21X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_18351_), .B(_19702__bF_buf4), .C(_19720_), .Y(_17347__17_) );
	OAI21X1 OAI21X1_4104 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf60), .Y(_19721_) );
	AOI21X1 AOI21X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_18405_), .B(_19702__bF_buf2), .C(_19721_), .Y(_17347__18_) );
	OAI21X1 OAI21X1_4105 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf59), .Y(_19722_) );
	AOI21X1 AOI21X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_18459_), .B(_19702__bF_buf0), .C(_19722_), .Y(_17347__19_) );
	OAI21X1 OAI21X1_4106 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf58), .Y(_19723_) );
	AOI21X1 AOI21X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_18513_), .B(_19702__bF_buf6), .C(_19723_), .Y(_17347__20_) );
	OAI21X1 OAI21X1_4107 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf57), .Y(_19724_) );
	AOI21X1 AOI21X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_18567_), .B(_19702__bF_buf4), .C(_19724_), .Y(_17347__21_) );
	OAI21X1 OAI21X1_4108 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf56), .Y(_19725_) );
	AOI21X1 AOI21X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_18621_), .B(_19702__bF_buf2), .C(_19725_), .Y(_17347__22_) );
	OAI21X1 OAI21X1_4109 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf55), .Y(_19726_) );
	AOI21X1 AOI21X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_18675_), .B(_19702__bF_buf0), .C(_19726_), .Y(_17347__23_) );
	OAI21X1 OAI21X1_4110 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf54), .Y(_19727_) );
	AOI21X1 AOI21X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_18729_), .B(_19702__bF_buf6), .C(_19727_), .Y(_17347__24_) );
	OAI21X1 OAI21X1_4111 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf53), .Y(_19728_) );
	AOI21X1 AOI21X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_18783_), .B(_19702__bF_buf4), .C(_19728_), .Y(_17347__25_) );
	OAI21X1 OAI21X1_4112 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf52), .Y(_19729_) );
	AOI21X1 AOI21X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_18837_), .B(_19702__bF_buf2), .C(_19729_), .Y(_17347__26_) );
	OAI21X1 OAI21X1_4113 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf51), .Y(_19730_) );
	AOI21X1 AOI21X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_18891_), .B(_19702__bF_buf0), .C(_19730_), .Y(_17347__27_) );
	OAI21X1 OAI21X1_4114 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf1), .B(_19702__bF_buf7), .C(_19153__bF_buf50), .Y(_19731_) );
	AOI21X1 AOI21X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_18945_), .B(_19702__bF_buf6), .C(_19731_), .Y(_17347__28_) );
	OAI21X1 OAI21X1_4115 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf1), .B(_19702__bF_buf5), .C(_19153__bF_buf49), .Y(_19732_) );
	AOI21X1 AOI21X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_18999_), .B(_19702__bF_buf4), .C(_19732_), .Y(_17347__29_) );
	OAI21X1 OAI21X1_4116 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf1), .B(_19702__bF_buf3), .C(_19153__bF_buf48), .Y(_19733_) );
	AOI21X1 AOI21X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_19053_), .B(_19702__bF_buf2), .C(_19733_), .Y(_17347__30_) );
	OAI21X1 OAI21X1_4117 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf1), .B(_19702__bF_buf1), .C(_19153__bF_buf47), .Y(_19734_) );
	AOI21X1 AOI21X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_19107_), .B(_19702__bF_buf0), .C(_19734_), .Y(_17347__31_) );
	NOR2X1 NOR2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_19254_), .B(_19666_), .Y(_19735_) );
	NAND2X1 NAND2X1_3558 ( .gnd(gnd), .vdd(vdd), .A(_19148_), .B(_19735_), .Y(_19736_) );
	OAI21X1 OAI21X1_4118 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf46), .Y(_19737_) );
	AOI21X1 AOI21X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_17453_), .B(_19736__bF_buf6), .C(_19737_), .Y(_17346__0_) );
	OAI21X1 OAI21X1_4119 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf45), .Y(_19738_) );
	AOI21X1 AOI21X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_17514_), .B(_19736__bF_buf4), .C(_19738_), .Y(_17346__1_) );
	OAI21X1 OAI21X1_4120 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf44), .Y(_19739_) );
	AOI21X1 AOI21X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_17568_), .B(_19736__bF_buf2), .C(_19739_), .Y(_17346__2_) );
	OAI21X1 OAI21X1_4121 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf43), .Y(_19740_) );
	AOI21X1 AOI21X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_17622_), .B(_19736__bF_buf0), .C(_19740_), .Y(_17346__3_) );
	OAI21X1 OAI21X1_4122 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf42), .Y(_19741_) );
	AOI21X1 AOI21X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_17676_), .B(_19736__bF_buf6), .C(_19741_), .Y(_17346__4_) );
	OAI21X1 OAI21X1_4123 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf41), .Y(_19742_) );
	AOI21X1 AOI21X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_17730_), .B(_19736__bF_buf4), .C(_19742_), .Y(_17346__5_) );
	OAI21X1 OAI21X1_4124 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf40), .Y(_19743_) );
	AOI21X1 AOI21X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_17784_), .B(_19736__bF_buf2), .C(_19743_), .Y(_17346__6_) );
	OAI21X1 OAI21X1_4125 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf39), .Y(_19744_) );
	AOI21X1 AOI21X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_17838_), .B(_19736__bF_buf0), .C(_19744_), .Y(_17346__7_) );
	OAI21X1 OAI21X1_4126 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf38), .Y(_19745_) );
	AOI21X1 AOI21X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_17892_), .B(_19736__bF_buf6), .C(_19745_), .Y(_17346__8_) );
	OAI21X1 OAI21X1_4127 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf37), .Y(_19746_) );
	AOI21X1 AOI21X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_17946_), .B(_19736__bF_buf4), .C(_19746_), .Y(_17346__9_) );
	OAI21X1 OAI21X1_4128 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf36), .Y(_19747_) );
	AOI21X1 AOI21X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_18000_), .B(_19736__bF_buf2), .C(_19747_), .Y(_17346__10_) );
	OAI21X1 OAI21X1_4129 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf35), .Y(_19748_) );
	AOI21X1 AOI21X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_18054_), .B(_19736__bF_buf0), .C(_19748_), .Y(_17346__11_) );
	OAI21X1 OAI21X1_4130 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf34), .Y(_19749_) );
	AOI21X1 AOI21X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_18108_), .B(_19736__bF_buf6), .C(_19749_), .Y(_17346__12_) );
	OAI21X1 OAI21X1_4131 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf33), .Y(_19750_) );
	AOI21X1 AOI21X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_18162_), .B(_19736__bF_buf4), .C(_19750_), .Y(_17346__13_) );
	OAI21X1 OAI21X1_4132 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf32), .Y(_19751_) );
	AOI21X1 AOI21X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_18216_), .B(_19736__bF_buf2), .C(_19751_), .Y(_17346__14_) );
	OAI21X1 OAI21X1_4133 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf31), .Y(_19752_) );
	AOI21X1 AOI21X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_18270_), .B(_19736__bF_buf0), .C(_19752_), .Y(_17346__15_) );
	OAI21X1 OAI21X1_4134 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf30), .Y(_19753_) );
	AOI21X1 AOI21X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_18324_), .B(_19736__bF_buf6), .C(_19753_), .Y(_17346__16_) );
	OAI21X1 OAI21X1_4135 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf29), .Y(_19754_) );
	AOI21X1 AOI21X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_18378_), .B(_19736__bF_buf4), .C(_19754_), .Y(_17346__17_) );
	OAI21X1 OAI21X1_4136 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf28), .Y(_19755_) );
	AOI21X1 AOI21X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_18432_), .B(_19736__bF_buf2), .C(_19755_), .Y(_17346__18_) );
	OAI21X1 OAI21X1_4137 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf27), .Y(_19756_) );
	AOI21X1 AOI21X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_18486_), .B(_19736__bF_buf0), .C(_19756_), .Y(_17346__19_) );
	OAI21X1 OAI21X1_4138 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf26), .Y(_19757_) );
	AOI21X1 AOI21X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_18540_), .B(_19736__bF_buf6), .C(_19757_), .Y(_17346__20_) );
	OAI21X1 OAI21X1_4139 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf25), .Y(_19758_) );
	AOI21X1 AOI21X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_18594_), .B(_19736__bF_buf4), .C(_19758_), .Y(_17346__21_) );
	OAI21X1 OAI21X1_4140 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf24), .Y(_19759_) );
	AOI21X1 AOI21X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_18648_), .B(_19736__bF_buf2), .C(_19759_), .Y(_17346__22_) );
	OAI21X1 OAI21X1_4141 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf23), .Y(_19760_) );
	AOI21X1 AOI21X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_18702_), .B(_19736__bF_buf0), .C(_19760_), .Y(_17346__23_) );
	OAI21X1 OAI21X1_4142 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf22), .Y(_19761_) );
	AOI21X1 AOI21X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_18756_), .B(_19736__bF_buf6), .C(_19761_), .Y(_17346__24_) );
	OAI21X1 OAI21X1_4143 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf21), .Y(_19762_) );
	AOI21X1 AOI21X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_18810_), .B(_19736__bF_buf4), .C(_19762_), .Y(_17346__25_) );
	OAI21X1 OAI21X1_4144 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf20), .Y(_19763_) );
	AOI21X1 AOI21X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_18864_), .B(_19736__bF_buf2), .C(_19763_), .Y(_17346__26_) );
	OAI21X1 OAI21X1_4145 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf19), .Y(_19764_) );
	AOI21X1 AOI21X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_18918_), .B(_19736__bF_buf0), .C(_19764_), .Y(_17346__27_) );
	OAI21X1 OAI21X1_4146 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf0), .B(_19736__bF_buf7), .C(_19153__bF_buf18), .Y(_19765_) );
	AOI21X1 AOI21X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_18972_), .B(_19736__bF_buf6), .C(_19765_), .Y(_17346__28_) );
	OAI21X1 OAI21X1_4147 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf0), .B(_19736__bF_buf5), .C(_19153__bF_buf17), .Y(_19766_) );
	AOI21X1 AOI21X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_19026_), .B(_19736__bF_buf4), .C(_19766_), .Y(_17346__29_) );
	OAI21X1 OAI21X1_4148 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf0), .B(_19736__bF_buf3), .C(_19153__bF_buf16), .Y(_19767_) );
	AOI21X1 AOI21X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_19080_), .B(_19736__bF_buf2), .C(_19767_), .Y(_17346__30_) );
	OAI21X1 OAI21X1_4149 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf0), .B(_19736__bF_buf1), .C(_19153__bF_buf15), .Y(_19768_) );
	AOI21X1 AOI21X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_19134_), .B(_19736__bF_buf0), .C(_19768_), .Y(_17346__31_) );
	NAND3X1 NAND3X1_3737 ( .gnd(gnd), .vdd(vdd), .A(_19496_), .B(_19325_), .C(_19430_), .Y(_19769_) );
	OAI21X1 OAI21X1_4150 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf14), .Y(_19770_) );
	AOI21X1 AOI21X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_17452_), .B(_19769__bF_buf6), .C(_19770_), .Y(_17345__0_) );
	OAI21X1 OAI21X1_4151 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf13), .Y(_19771_) );
	AOI21X1 AOI21X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_17513_), .B(_19769__bF_buf4), .C(_19771_), .Y(_17345__1_) );
	OAI21X1 OAI21X1_4152 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf12), .Y(_19772_) );
	AOI21X1 AOI21X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_17567_), .B(_19769__bF_buf2), .C(_19772_), .Y(_17345__2_) );
	OAI21X1 OAI21X1_4153 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf11), .Y(_19773_) );
	AOI21X1 AOI21X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_17621_), .B(_19769__bF_buf0), .C(_19773_), .Y(_17345__3_) );
	OAI21X1 OAI21X1_4154 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf10), .Y(_19774_) );
	AOI21X1 AOI21X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_17675_), .B(_19769__bF_buf6), .C(_19774_), .Y(_17345__4_) );
	OAI21X1 OAI21X1_4155 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf9), .Y(_19775_) );
	AOI21X1 AOI21X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_17729_), .B(_19769__bF_buf4), .C(_19775_), .Y(_17345__5_) );
	OAI21X1 OAI21X1_4156 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf8), .Y(_19776_) );
	AOI21X1 AOI21X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_17783_), .B(_19769__bF_buf2), .C(_19776_), .Y(_17345__6_) );
	OAI21X1 OAI21X1_4157 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf7), .Y(_19777_) );
	AOI21X1 AOI21X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_17837_), .B(_19769__bF_buf0), .C(_19777_), .Y(_17345__7_) );
	OAI21X1 OAI21X1_4158 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf6), .Y(_19778_) );
	AOI21X1 AOI21X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_17891_), .B(_19769__bF_buf6), .C(_19778_), .Y(_17345__8_) );
	OAI21X1 OAI21X1_4159 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf5), .Y(_19779_) );
	AOI21X1 AOI21X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_17945_), .B(_19769__bF_buf4), .C(_19779_), .Y(_17345__9_) );
	OAI21X1 OAI21X1_4160 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf4), .Y(_19780_) );
	AOI21X1 AOI21X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_17999_), .B(_19769__bF_buf2), .C(_19780_), .Y(_17345__10_) );
	OAI21X1 OAI21X1_4161 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf3), .Y(_19781_) );
	AOI21X1 AOI21X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_18053_), .B(_19769__bF_buf0), .C(_19781_), .Y(_17345__11_) );
	OAI21X1 OAI21X1_4162 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf2), .Y(_19782_) );
	AOI21X1 AOI21X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_18107_), .B(_19769__bF_buf6), .C(_19782_), .Y(_17345__12_) );
	OAI21X1 OAI21X1_4163 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf1), .Y(_19783_) );
	AOI21X1 AOI21X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_18161_), .B(_19769__bF_buf4), .C(_19783_), .Y(_17345__13_) );
	OAI21X1 OAI21X1_4164 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf0), .Y(_19784_) );
	AOI21X1 AOI21X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_18215_), .B(_19769__bF_buf2), .C(_19784_), .Y(_17345__14_) );
	OAI21X1 OAI21X1_4165 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf98), .Y(_19785_) );
	AOI21X1 AOI21X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_18269_), .B(_19769__bF_buf0), .C(_19785_), .Y(_17345__15_) );
	OAI21X1 OAI21X1_4166 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf97), .Y(_19786_) );
	AOI21X1 AOI21X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_18323_), .B(_19769__bF_buf6), .C(_19786_), .Y(_17345__16_) );
	OAI21X1 OAI21X1_4167 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf96), .Y(_19787_) );
	AOI21X1 AOI21X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_18377_), .B(_19769__bF_buf4), .C(_19787_), .Y(_17345__17_) );
	OAI21X1 OAI21X1_4168 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf95), .Y(_19788_) );
	AOI21X1 AOI21X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_18431_), .B(_19769__bF_buf2), .C(_19788_), .Y(_17345__18_) );
	OAI21X1 OAI21X1_4169 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf94), .Y(_19789_) );
	AOI21X1 AOI21X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_18485_), .B(_19769__bF_buf0), .C(_19789_), .Y(_17345__19_) );
	OAI21X1 OAI21X1_4170 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf93), .Y(_19790_) );
	AOI21X1 AOI21X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_18539_), .B(_19769__bF_buf6), .C(_19790_), .Y(_17345__20_) );
	OAI21X1 OAI21X1_4171 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf92), .Y(_19791_) );
	AOI21X1 AOI21X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_18593_), .B(_19769__bF_buf4), .C(_19791_), .Y(_17345__21_) );
	OAI21X1 OAI21X1_4172 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf91), .Y(_19792_) );
	AOI21X1 AOI21X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_18647_), .B(_19769__bF_buf2), .C(_19792_), .Y(_17345__22_) );
	OAI21X1 OAI21X1_4173 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf90), .Y(_19793_) );
	AOI21X1 AOI21X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_18701_), .B(_19769__bF_buf0), .C(_19793_), .Y(_17345__23_) );
	OAI21X1 OAI21X1_4174 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf89), .Y(_19794_) );
	AOI21X1 AOI21X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_18755_), .B(_19769__bF_buf6), .C(_19794_), .Y(_17345__24_) );
	OAI21X1 OAI21X1_4175 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf88), .Y(_19795_) );
	AOI21X1 AOI21X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_18809_), .B(_19769__bF_buf4), .C(_19795_), .Y(_17345__25_) );
	OAI21X1 OAI21X1_4176 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf87), .Y(_19796_) );
	AOI21X1 AOI21X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_18863_), .B(_19769__bF_buf2), .C(_19796_), .Y(_17345__26_) );
	OAI21X1 OAI21X1_4177 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf86), .Y(_19797_) );
	AOI21X1 AOI21X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_18917_), .B(_19769__bF_buf0), .C(_19797_), .Y(_17345__27_) );
	OAI21X1 OAI21X1_4178 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_19769__bF_buf7), .C(_19153__bF_buf85), .Y(_19798_) );
	AOI21X1 AOI21X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_18971_), .B(_19769__bF_buf6), .C(_19798_), .Y(_17345__28_) );
	OAI21X1 OAI21X1_4179 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_19769__bF_buf5), .C(_19153__bF_buf84), .Y(_19799_) );
	AOI21X1 AOI21X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_19025_), .B(_19769__bF_buf4), .C(_19799_), .Y(_17345__29_) );
	OAI21X1 OAI21X1_4180 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_19769__bF_buf3), .C(_19153__bF_buf83), .Y(_19800_) );
	AOI21X1 AOI21X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_19079_), .B(_19769__bF_buf2), .C(_19800_), .Y(_17345__30_) );
	OAI21X1 OAI21X1_4181 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_19769__bF_buf1), .C(_19153__bF_buf82), .Y(_19801_) );
	AOI21X1 AOI21X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_19133_), .B(_19769__bF_buf0), .C(_19801_), .Y(_17345__31_) );
	INVX1 INVX1_2881 ( .gnd(gnd), .vdd(vdd), .A(registers_writeEnable), .Y(_19802_) );
	NOR2X1 NOR2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(instructionFrame_writeSelect_out_4_), .B(_19802_), .Y(_19803_) );
	NAND2X1 NAND2X1_3559 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19151_), .Y(_19804_) );
	OAI21X1 OAI21X1_4182 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf81), .Y(_19805_) );
	AOI21X1 AOI21X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_17441_), .B(_19804__bF_buf6), .C(_19805_), .Y(_17344__0_) );
	OAI21X1 OAI21X1_4183 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf80), .Y(_19806_) );
	AOI21X1 AOI21X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_17505_), .B(_19804__bF_buf4), .C(_19806_), .Y(_17344__1_) );
	OAI21X1 OAI21X1_4184 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf79), .Y(_19807_) );
	AOI21X1 AOI21X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_17559_), .B(_19804__bF_buf2), .C(_19807_), .Y(_17344__2_) );
	OAI21X1 OAI21X1_4185 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf78), .Y(_19808_) );
	AOI21X1 AOI21X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_17613_), .B(_19804__bF_buf0), .C(_19808_), .Y(_17344__3_) );
	OAI21X1 OAI21X1_4186 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf77), .Y(_19809_) );
	AOI21X1 AOI21X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_17667_), .B(_19804__bF_buf6), .C(_19809_), .Y(_17344__4_) );
	OAI21X1 OAI21X1_4187 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf76), .Y(_19810_) );
	AOI21X1 AOI21X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_17721_), .B(_19804__bF_buf4), .C(_19810_), .Y(_17344__5_) );
	OAI21X1 OAI21X1_4188 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf75), .Y(_19811_) );
	AOI21X1 AOI21X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_17775_), .B(_19804__bF_buf2), .C(_19811_), .Y(_17344__6_) );
	OAI21X1 OAI21X1_4189 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf74), .Y(_19812_) );
	AOI21X1 AOI21X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_17829_), .B(_19804__bF_buf0), .C(_19812_), .Y(_17344__7_) );
	OAI21X1 OAI21X1_4190 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf73), .Y(_19813_) );
	AOI21X1 AOI21X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_17883_), .B(_19804__bF_buf6), .C(_19813_), .Y(_17344__8_) );
	OAI21X1 OAI21X1_4191 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf72), .Y(_19814_) );
	AOI21X1 AOI21X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_17937_), .B(_19804__bF_buf4), .C(_19814_), .Y(_17344__9_) );
	OAI21X1 OAI21X1_4192 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf71), .Y(_19815_) );
	AOI21X1 AOI21X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_17991_), .B(_19804__bF_buf2), .C(_19815_), .Y(_17344__10_) );
	OAI21X1 OAI21X1_4193 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf70), .Y(_19816_) );
	AOI21X1 AOI21X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_18045_), .B(_19804__bF_buf0), .C(_19816_), .Y(_17344__11_) );
	OAI21X1 OAI21X1_4194 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf69), .Y(_19817_) );
	AOI21X1 AOI21X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_18099_), .B(_19804__bF_buf6), .C(_19817_), .Y(_17344__12_) );
	OAI21X1 OAI21X1_4195 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf68), .Y(_19818_) );
	AOI21X1 AOI21X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_18153_), .B(_19804__bF_buf4), .C(_19818_), .Y(_17344__13_) );
	OAI21X1 OAI21X1_4196 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf67), .Y(_19819_) );
	AOI21X1 AOI21X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_18207_), .B(_19804__bF_buf2), .C(_19819_), .Y(_17344__14_) );
	OAI21X1 OAI21X1_4197 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf66), .Y(_19820_) );
	AOI21X1 AOI21X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_18261_), .B(_19804__bF_buf0), .C(_19820_), .Y(_17344__15_) );
	OAI21X1 OAI21X1_4198 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf65), .Y(_19821_) );
	AOI21X1 AOI21X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_18315_), .B(_19804__bF_buf6), .C(_19821_), .Y(_17344__16_) );
	OAI21X1 OAI21X1_4199 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf64), .Y(_19822_) );
	AOI21X1 AOI21X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_18369_), .B(_19804__bF_buf4), .C(_19822_), .Y(_17344__17_) );
	OAI21X1 OAI21X1_4200 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf63), .Y(_19823_) );
	AOI21X1 AOI21X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_18423_), .B(_19804__bF_buf2), .C(_19823_), .Y(_17344__18_) );
	OAI21X1 OAI21X1_4201 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf62), .Y(_19824_) );
	AOI21X1 AOI21X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_18477_), .B(_19804__bF_buf0), .C(_19824_), .Y(_17344__19_) );
	OAI21X1 OAI21X1_4202 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf61), .Y(_19825_) );
	AOI21X1 AOI21X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_18531_), .B(_19804__bF_buf6), .C(_19825_), .Y(_17344__20_) );
	OAI21X1 OAI21X1_4203 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf60), .Y(_19826_) );
	AOI21X1 AOI21X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_18585_), .B(_19804__bF_buf4), .C(_19826_), .Y(_17344__21_) );
	OAI21X1 OAI21X1_4204 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf59), .Y(_19827_) );
	AOI21X1 AOI21X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_18639_), .B(_19804__bF_buf2), .C(_19827_), .Y(_17344__22_) );
	OAI21X1 OAI21X1_4205 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf58), .Y(_19828_) );
	AOI21X1 AOI21X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_18693_), .B(_19804__bF_buf0), .C(_19828_), .Y(_17344__23_) );
	OAI21X1 OAI21X1_4206 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf57), .Y(_19829_) );
	AOI21X1 AOI21X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_18747_), .B(_19804__bF_buf6), .C(_19829_), .Y(_17344__24_) );
	OAI21X1 OAI21X1_4207 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf56), .Y(_19830_) );
	AOI21X1 AOI21X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_18801_), .B(_19804__bF_buf4), .C(_19830_), .Y(_17344__25_) );
	OAI21X1 OAI21X1_4208 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf55), .Y(_19831_) );
	AOI21X1 AOI21X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_18855_), .B(_19804__bF_buf2), .C(_19831_), .Y(_17344__26_) );
	OAI21X1 OAI21X1_4209 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf54), .Y(_19832_) );
	AOI21X1 AOI21X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_18909_), .B(_19804__bF_buf0), .C(_19832_), .Y(_17344__27_) );
	OAI21X1 OAI21X1_4210 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf3), .B(_19804__bF_buf7), .C(_19153__bF_buf53), .Y(_19833_) );
	AOI21X1 AOI21X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_18963_), .B(_19804__bF_buf6), .C(_19833_), .Y(_17344__28_) );
	OAI21X1 OAI21X1_4211 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf3), .B(_19804__bF_buf5), .C(_19153__bF_buf52), .Y(_19834_) );
	AOI21X1 AOI21X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_19017_), .B(_19804__bF_buf4), .C(_19834_), .Y(_17344__29_) );
	OAI21X1 OAI21X1_4212 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf3), .B(_19804__bF_buf3), .C(_19153__bF_buf51), .Y(_19835_) );
	AOI21X1 AOI21X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_19071_), .B(_19804__bF_buf2), .C(_19835_), .Y(_17344__30_) );
	OAI21X1 OAI21X1_4213 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf3), .B(_19804__bF_buf1), .C(_19153__bF_buf50), .Y(_19836_) );
	AOI21X1 AOI21X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_19125_), .B(_19804__bF_buf0), .C(_19836_), .Y(_17344__31_) );
	NAND2X1 NAND2X1_3560 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19219_), .Y(_19837_) );
	OAI21X1 OAI21X1_4214 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf49), .Y(_19838_) );
	AOI21X1 AOI21X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_17396_), .B(_19837__bF_buf6), .C(_19838_), .Y(_17343__0_) );
	OAI21X1 OAI21X1_4215 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf48), .Y(_19839_) );
	AOI21X1 AOI21X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_17482_), .B(_19837__bF_buf4), .C(_19839_), .Y(_17343__1_) );
	OAI21X1 OAI21X1_4216 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf47), .Y(_19840_) );
	AOI21X1 AOI21X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_17536_), .B(_19837__bF_buf2), .C(_19840_), .Y(_17343__2_) );
	OAI21X1 OAI21X1_4217 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf46), .Y(_19841_) );
	AOI21X1 AOI21X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_17590_), .B(_19837__bF_buf0), .C(_19841_), .Y(_17343__3_) );
	OAI21X1 OAI21X1_4218 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf45), .Y(_19842_) );
	AOI21X1 AOI21X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_17644_), .B(_19837__bF_buf6), .C(_19842_), .Y(_17343__4_) );
	OAI21X1 OAI21X1_4219 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf44), .Y(_19843_) );
	AOI21X1 AOI21X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_17698_), .B(_19837__bF_buf4), .C(_19843_), .Y(_17343__5_) );
	OAI21X1 OAI21X1_4220 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf43), .Y(_19844_) );
	AOI21X1 AOI21X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_17752_), .B(_19837__bF_buf2), .C(_19844_), .Y(_17343__6_) );
	OAI21X1 OAI21X1_4221 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf42), .Y(_19845_) );
	AOI21X1 AOI21X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_17806_), .B(_19837__bF_buf0), .C(_19845_), .Y(_17343__7_) );
	OAI21X1 OAI21X1_4222 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf41), .Y(_19846_) );
	AOI21X1 AOI21X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_17860_), .B(_19837__bF_buf6), .C(_19846_), .Y(_17343__8_) );
	OAI21X1 OAI21X1_4223 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf40), .Y(_19847_) );
	AOI21X1 AOI21X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_17914_), .B(_19837__bF_buf4), .C(_19847_), .Y(_17343__9_) );
	OAI21X1 OAI21X1_4224 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf39), .Y(_19848_) );
	AOI21X1 AOI21X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_17968_), .B(_19837__bF_buf2), .C(_19848_), .Y(_17343__10_) );
	OAI21X1 OAI21X1_4225 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf38), .Y(_19849_) );
	AOI21X1 AOI21X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_18022_), .B(_19837__bF_buf0), .C(_19849_), .Y(_17343__11_) );
	OAI21X1 OAI21X1_4226 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf37), .Y(_19850_) );
	AOI21X1 AOI21X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_18076_), .B(_19837__bF_buf6), .C(_19850_), .Y(_17343__12_) );
	OAI21X1 OAI21X1_4227 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf36), .Y(_19851_) );
	AOI21X1 AOI21X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_18130_), .B(_19837__bF_buf4), .C(_19851_), .Y(_17343__13_) );
	OAI21X1 OAI21X1_4228 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf35), .Y(_19852_) );
	AOI21X1 AOI21X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_18184_), .B(_19837__bF_buf2), .C(_19852_), .Y(_17343__14_) );
	OAI21X1 OAI21X1_4229 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf34), .Y(_19853_) );
	AOI21X1 AOI21X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_18238_), .B(_19837__bF_buf0), .C(_19853_), .Y(_17343__15_) );
	OAI21X1 OAI21X1_4230 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf33), .Y(_19854_) );
	AOI21X1 AOI21X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_18292_), .B(_19837__bF_buf6), .C(_19854_), .Y(_17343__16_) );
	OAI21X1 OAI21X1_4231 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf32), .Y(_19855_) );
	AOI21X1 AOI21X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_18346_), .B(_19837__bF_buf4), .C(_19855_), .Y(_17343__17_) );
	OAI21X1 OAI21X1_4232 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf31), .Y(_19856_) );
	AOI21X1 AOI21X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_18400_), .B(_19837__bF_buf2), .C(_19856_), .Y(_17343__18_) );
	OAI21X1 OAI21X1_4233 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf30), .Y(_19857_) );
	AOI21X1 AOI21X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_18454_), .B(_19837__bF_buf0), .C(_19857_), .Y(_17343__19_) );
	OAI21X1 OAI21X1_4234 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf29), .Y(_19858_) );
	AOI21X1 AOI21X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_18508_), .B(_19837__bF_buf6), .C(_19858_), .Y(_17343__20_) );
	OAI21X1 OAI21X1_4235 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf28), .Y(_19859_) );
	AOI21X1 AOI21X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_18562_), .B(_19837__bF_buf4), .C(_19859_), .Y(_17343__21_) );
	OAI21X1 OAI21X1_4236 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf27), .Y(_19860_) );
	AOI21X1 AOI21X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_18616_), .B(_19837__bF_buf2), .C(_19860_), .Y(_17343__22_) );
	OAI21X1 OAI21X1_4237 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf26), .Y(_19861_) );
	AOI21X1 AOI21X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_18670_), .B(_19837__bF_buf0), .C(_19861_), .Y(_17343__23_) );
	OAI21X1 OAI21X1_4238 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf25), .Y(_19862_) );
	AOI21X1 AOI21X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_18724_), .B(_19837__bF_buf6), .C(_19862_), .Y(_17343__24_) );
	OAI21X1 OAI21X1_4239 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf24), .Y(_19863_) );
	AOI21X1 AOI21X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_18778_), .B(_19837__bF_buf4), .C(_19863_), .Y(_17343__25_) );
	OAI21X1 OAI21X1_4240 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf23), .Y(_19864_) );
	AOI21X1 AOI21X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_18832_), .B(_19837__bF_buf2), .C(_19864_), .Y(_17343__26_) );
	OAI21X1 OAI21X1_4241 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf22), .Y(_19865_) );
	AOI21X1 AOI21X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_18886_), .B(_19837__bF_buf0), .C(_19865_), .Y(_17343__27_) );
	OAI21X1 OAI21X1_4242 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf2), .B(_19837__bF_buf7), .C(_19153__bF_buf21), .Y(_19866_) );
	AOI21X1 AOI21X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_18940_), .B(_19837__bF_buf6), .C(_19866_), .Y(_17343__28_) );
	OAI21X1 OAI21X1_4243 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf2), .B(_19837__bF_buf5), .C(_19153__bF_buf20), .Y(_19867_) );
	AOI21X1 AOI21X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_18994_), .B(_19837__bF_buf4), .C(_19867_), .Y(_17343__29_) );
	OAI21X1 OAI21X1_4244 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf2), .B(_19837__bF_buf3), .C(_19153__bF_buf19), .Y(_19868_) );
	AOI21X1 AOI21X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_19048_), .B(_19837__bF_buf2), .C(_19868_), .Y(_17343__30_) );
	OAI21X1 OAI21X1_4245 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf2), .B(_19837__bF_buf1), .C(_19153__bF_buf18), .Y(_19869_) );
	AOI21X1 AOI21X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_19102_), .B(_19837__bF_buf0), .C(_19869_), .Y(_17343__31_) );
	NAND2X1 NAND2X1_3561 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19255_), .Y(_19870_) );
	OAI21X1 OAI21X1_4246 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf17), .Y(_19871_) );
	AOI21X1 AOI21X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_17397_), .B(_19870__bF_buf6), .C(_19871_), .Y(_17342__0_) );
	OAI21X1 OAI21X1_4247 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf16), .Y(_19872_) );
	AOI21X1 AOI21X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_17483_), .B(_19870__bF_buf4), .C(_19872_), .Y(_17342__1_) );
	OAI21X1 OAI21X1_4248 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf15), .Y(_19873_) );
	AOI21X1 AOI21X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_17537_), .B(_19870__bF_buf2), .C(_19873_), .Y(_17342__2_) );
	OAI21X1 OAI21X1_4249 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf14), .Y(_19874_) );
	AOI21X1 AOI21X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_17591_), .B(_19870__bF_buf0), .C(_19874_), .Y(_17342__3_) );
	OAI21X1 OAI21X1_4250 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf13), .Y(_19875_) );
	AOI21X1 AOI21X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_17645_), .B(_19870__bF_buf6), .C(_19875_), .Y(_17342__4_) );
	OAI21X1 OAI21X1_4251 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf12), .Y(_19876_) );
	AOI21X1 AOI21X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_17699_), .B(_19870__bF_buf4), .C(_19876_), .Y(_17342__5_) );
	OAI21X1 OAI21X1_4252 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf11), .Y(_19877_) );
	AOI21X1 AOI21X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_17753_), .B(_19870__bF_buf2), .C(_19877_), .Y(_17342__6_) );
	OAI21X1 OAI21X1_4253 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf10), .Y(_19878_) );
	AOI21X1 AOI21X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_17807_), .B(_19870__bF_buf0), .C(_19878_), .Y(_17342__7_) );
	OAI21X1 OAI21X1_4254 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf9), .Y(_19879_) );
	AOI21X1 AOI21X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_17861_), .B(_19870__bF_buf6), .C(_19879_), .Y(_17342__8_) );
	OAI21X1 OAI21X1_4255 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf8), .Y(_19880_) );
	AOI21X1 AOI21X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_17915_), .B(_19870__bF_buf4), .C(_19880_), .Y(_17342__9_) );
	OAI21X1 OAI21X1_4256 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf7), .Y(_19881_) );
	AOI21X1 AOI21X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_17969_), .B(_19870__bF_buf2), .C(_19881_), .Y(_17342__10_) );
	OAI21X1 OAI21X1_4257 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf6), .Y(_19882_) );
	AOI21X1 AOI21X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_18023_), .B(_19870__bF_buf0), .C(_19882_), .Y(_17342__11_) );
	OAI21X1 OAI21X1_4258 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf5), .Y(_19883_) );
	AOI21X1 AOI21X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_18077_), .B(_19870__bF_buf6), .C(_19883_), .Y(_17342__12_) );
	OAI21X1 OAI21X1_4259 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf4), .Y(_19884_) );
	AOI21X1 AOI21X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_18131_), .B(_19870__bF_buf4), .C(_19884_), .Y(_17342__13_) );
	OAI21X1 OAI21X1_4260 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf3), .Y(_19885_) );
	AOI21X1 AOI21X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_18185_), .B(_19870__bF_buf2), .C(_19885_), .Y(_17342__14_) );
	OAI21X1 OAI21X1_4261 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf2), .Y(_19886_) );
	AOI21X1 AOI21X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_18239_), .B(_19870__bF_buf0), .C(_19886_), .Y(_17342__15_) );
	OAI21X1 OAI21X1_4262 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf1), .Y(_19887_) );
	AOI21X1 AOI21X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_18293_), .B(_19870__bF_buf6), .C(_19887_), .Y(_17342__16_) );
	OAI21X1 OAI21X1_4263 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf0), .Y(_19888_) );
	AOI21X1 AOI21X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_18347_), .B(_19870__bF_buf4), .C(_19888_), .Y(_17342__17_) );
	OAI21X1 OAI21X1_4264 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf98), .Y(_19889_) );
	AOI21X1 AOI21X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_18401_), .B(_19870__bF_buf2), .C(_19889_), .Y(_17342__18_) );
	OAI21X1 OAI21X1_4265 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf97), .Y(_19890_) );
	AOI21X1 AOI21X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_18455_), .B(_19870__bF_buf0), .C(_19890_), .Y(_17342__19_) );
	OAI21X1 OAI21X1_4266 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf96), .Y(_19891_) );
	AOI21X1 AOI21X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_18509_), .B(_19870__bF_buf6), .C(_19891_), .Y(_17342__20_) );
	OAI21X1 OAI21X1_4267 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf95), .Y(_19892_) );
	AOI21X1 AOI21X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_18563_), .B(_19870__bF_buf4), .C(_19892_), .Y(_17342__21_) );
	OAI21X1 OAI21X1_4268 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf94), .Y(_19893_) );
	AOI21X1 AOI21X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_18617_), .B(_19870__bF_buf2), .C(_19893_), .Y(_17342__22_) );
	OAI21X1 OAI21X1_4269 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf93), .Y(_19894_) );
	AOI21X1 AOI21X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_18671_), .B(_19870__bF_buf0), .C(_19894_), .Y(_17342__23_) );
	OAI21X1 OAI21X1_4270 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf92), .Y(_19895_) );
	AOI21X1 AOI21X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_18725_), .B(_19870__bF_buf6), .C(_19895_), .Y(_17342__24_) );
	OAI21X1 OAI21X1_4271 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf91), .Y(_19896_) );
	AOI21X1 AOI21X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_18779_), .B(_19870__bF_buf4), .C(_19896_), .Y(_17342__25_) );
	OAI21X1 OAI21X1_4272 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf90), .Y(_19897_) );
	AOI21X1 AOI21X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_18833_), .B(_19870__bF_buf2), .C(_19897_), .Y(_17342__26_) );
	OAI21X1 OAI21X1_4273 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf89), .Y(_19898_) );
	AOI21X1 AOI21X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_18887_), .B(_19870__bF_buf0), .C(_19898_), .Y(_17342__27_) );
	OAI21X1 OAI21X1_4274 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf1), .B(_19870__bF_buf7), .C(_19153__bF_buf88), .Y(_19899_) );
	AOI21X1 AOI21X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_18941_), .B(_19870__bF_buf6), .C(_19899_), .Y(_17342__28_) );
	OAI21X1 OAI21X1_4275 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf1), .B(_19870__bF_buf5), .C(_19153__bF_buf87), .Y(_19900_) );
	AOI21X1 AOI21X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_18995_), .B(_19870__bF_buf4), .C(_19900_), .Y(_17342__29_) );
	OAI21X1 OAI21X1_4276 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf1), .B(_19870__bF_buf3), .C(_19153__bF_buf86), .Y(_19901_) );
	AOI21X1 AOI21X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_19049_), .B(_19870__bF_buf2), .C(_19901_), .Y(_17342__30_) );
	OAI21X1 OAI21X1_4277 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf1), .B(_19870__bF_buf1), .C(_19153__bF_buf85), .Y(_19902_) );
	AOI21X1 AOI21X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_19103_), .B(_19870__bF_buf0), .C(_19902_), .Y(_17342__31_) );
	INVX1 INVX1_2882 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_0_), .Y(_19903_) );
	NAND2X1 NAND2X1_3562 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19291_), .Y(_19904_) );
	OAI21X1 OAI21X1_4278 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf84), .Y(_19905_) );
	AOI21X1 AOI21X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_19903_), .B(_19904__bF_buf6), .C(_19905_), .Y(_17341__0_) );
	INVX1 INVX1_2883 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_1_), .Y(_19906_) );
	OAI21X1 OAI21X1_4279 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf83), .Y(_19907_) );
	AOI21X1 AOI21X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_19906_), .B(_19904__bF_buf4), .C(_19907_), .Y(_17341__1_) );
	INVX1 INVX1_2884 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_2_), .Y(_19908_) );
	OAI21X1 OAI21X1_4280 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf82), .Y(_19909_) );
	AOI21X1 AOI21X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_19908_), .B(_19904__bF_buf2), .C(_19909_), .Y(_17341__2_) );
	INVX1 INVX1_2885 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_3_), .Y(_19910_) );
	OAI21X1 OAI21X1_4281 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf81), .Y(_19911_) );
	AOI21X1 AOI21X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_19910_), .B(_19904__bF_buf0), .C(_19911_), .Y(_17341__3_) );
	INVX1 INVX1_2886 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_4_), .Y(_19912_) );
	OAI21X1 OAI21X1_4282 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf80), .Y(_19913_) );
	AOI21X1 AOI21X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_19912_), .B(_19904__bF_buf6), .C(_19913_), .Y(_17341__4_) );
	INVX1 INVX1_2887 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_5_), .Y(_19914_) );
	OAI21X1 OAI21X1_4283 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf79), .Y(_19915_) );
	AOI21X1 AOI21X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_19914_), .B(_19904__bF_buf4), .C(_19915_), .Y(_17341__5_) );
	INVX1 INVX1_2888 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_6_), .Y(_19916_) );
	OAI21X1 OAI21X1_4284 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf78), .Y(_19917_) );
	AOI21X1 AOI21X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_19916_), .B(_19904__bF_buf2), .C(_19917_), .Y(_17341__6_) );
	INVX1 INVX1_2889 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_7_), .Y(_19918_) );
	OAI21X1 OAI21X1_4285 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf77), .Y(_19919_) );
	AOI21X1 AOI21X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_19918_), .B(_19904__bF_buf0), .C(_19919_), .Y(_17341__7_) );
	INVX1 INVX1_2890 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_8_), .Y(_19920_) );
	OAI21X1 OAI21X1_4286 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf76), .Y(_19921_) );
	AOI21X1 AOI21X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_19920_), .B(_19904__bF_buf6), .C(_19921_), .Y(_17341__8_) );
	INVX1 INVX1_2891 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_9_), .Y(_19922_) );
	OAI21X1 OAI21X1_4287 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf75), .Y(_19923_) );
	AOI21X1 AOI21X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_19922_), .B(_19904__bF_buf4), .C(_19923_), .Y(_17341__9_) );
	INVX1 INVX1_2892 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_10_), .Y(_19924_) );
	OAI21X1 OAI21X1_4288 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf74), .Y(_19925_) );
	AOI21X1 AOI21X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_19924_), .B(_19904__bF_buf2), .C(_19925_), .Y(_17341__10_) );
	INVX1 INVX1_2893 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_11_), .Y(_19926_) );
	OAI21X1 OAI21X1_4289 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf73), .Y(_19927_) );
	AOI21X1 AOI21X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_19926_), .B(_19904__bF_buf0), .C(_19927_), .Y(_17341__11_) );
	INVX1 INVX1_2894 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_12_), .Y(_19928_) );
	OAI21X1 OAI21X1_4290 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf72), .Y(_19929_) );
	AOI21X1 AOI21X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_19928_), .B(_19904__bF_buf6), .C(_19929_), .Y(_17341__12_) );
	INVX1 INVX1_2895 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_13_), .Y(_19930_) );
	OAI21X1 OAI21X1_4291 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf71), .Y(_19931_) );
	AOI21X1 AOI21X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_19930_), .B(_19904__bF_buf4), .C(_19931_), .Y(_17341__13_) );
	INVX1 INVX1_2896 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_14_), .Y(_19932_) );
	OAI21X1 OAI21X1_4292 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf70), .Y(_19933_) );
	AOI21X1 AOI21X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_19932_), .B(_19904__bF_buf2), .C(_19933_), .Y(_17341__14_) );
	INVX1 INVX1_2897 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_15_), .Y(_19934_) );
	OAI21X1 OAI21X1_4293 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf69), .Y(_19935_) );
	AOI21X1 AOI21X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_19934_), .B(_19904__bF_buf0), .C(_19935_), .Y(_17341__15_) );
	INVX1 INVX1_2898 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_16_), .Y(_19936_) );
	OAI21X1 OAI21X1_4294 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf68), .Y(_19937_) );
	AOI21X1 AOI21X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_19936_), .B(_19904__bF_buf6), .C(_19937_), .Y(_17341__16_) );
	INVX1 INVX1_2899 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_17_), .Y(_19938_) );
	OAI21X1 OAI21X1_4295 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf67), .Y(_19939_) );
	AOI21X1 AOI21X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_19938_), .B(_19904__bF_buf4), .C(_19939_), .Y(_17341__17_) );
	INVX1 INVX1_2900 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_18_), .Y(_19940_) );
	OAI21X1 OAI21X1_4296 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf66), .Y(_19941_) );
	AOI21X1 AOI21X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_19940_), .B(_19904__bF_buf2), .C(_19941_), .Y(_17341__18_) );
	INVX1 INVX1_2901 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_19_), .Y(_19942_) );
	OAI21X1 OAI21X1_4297 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf65), .Y(_19943_) );
	AOI21X1 AOI21X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_19942_), .B(_19904__bF_buf0), .C(_19943_), .Y(_17341__19_) );
	INVX1 INVX1_2902 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_20_), .Y(_19944_) );
	OAI21X1 OAI21X1_4298 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf64), .Y(_19945_) );
	AOI21X1 AOI21X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_19944_), .B(_19904__bF_buf6), .C(_19945_), .Y(_17341__20_) );
	INVX1 INVX1_2903 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_21_), .Y(_19946_) );
	OAI21X1 OAI21X1_4299 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf63), .Y(_19947_) );
	AOI21X1 AOI21X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_19946_), .B(_19904__bF_buf4), .C(_19947_), .Y(_17341__21_) );
	INVX1 INVX1_2904 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_22_), .Y(_19948_) );
	OAI21X1 OAI21X1_4300 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf62), .Y(_19949_) );
	AOI21X1 AOI21X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_19948_), .B(_19904__bF_buf2), .C(_19949_), .Y(_17341__22_) );
	INVX1 INVX1_2905 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_23_), .Y(_19950_) );
	OAI21X1 OAI21X1_4301 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf61), .Y(_19951_) );
	AOI21X1 AOI21X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_19950_), .B(_19904__bF_buf0), .C(_19951_), .Y(_17341__23_) );
	INVX1 INVX1_2906 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_24_), .Y(_19952_) );
	OAI21X1 OAI21X1_4302 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf60), .Y(_19953_) );
	AOI21X1 AOI21X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_19952_), .B(_19904__bF_buf6), .C(_19953_), .Y(_17341__24_) );
	INVX1 INVX1_2907 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_25_), .Y(_19954_) );
	OAI21X1 OAI21X1_4303 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf59), .Y(_19955_) );
	AOI21X1 AOI21X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_19954_), .B(_19904__bF_buf4), .C(_19955_), .Y(_17341__25_) );
	INVX1 INVX1_2908 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_26_), .Y(_19956_) );
	OAI21X1 OAI21X1_4304 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf58), .Y(_19957_) );
	AOI21X1 AOI21X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_19956_), .B(_19904__bF_buf2), .C(_19957_), .Y(_17341__26_) );
	INVX1 INVX1_2909 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_27_), .Y(_19958_) );
	OAI21X1 OAI21X1_4305 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf57), .Y(_19959_) );
	AOI21X1 AOI21X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_19958_), .B(_19904__bF_buf0), .C(_19959_), .Y(_17341__27_) );
	INVX1 INVX1_2910 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_28_), .Y(_19960_) );
	OAI21X1 OAI21X1_4306 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf0), .B(_19904__bF_buf7), .C(_19153__bF_buf56), .Y(_19961_) );
	AOI21X1 AOI21X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_19960_), .B(_19904__bF_buf6), .C(_19961_), .Y(_17341__28_) );
	INVX1 INVX1_2911 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_29_), .Y(_19962_) );
	OAI21X1 OAI21X1_4307 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf0), .B(_19904__bF_buf5), .C(_19153__bF_buf55), .Y(_19963_) );
	AOI21X1 AOI21X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_19962_), .B(_19904__bF_buf4), .C(_19963_), .Y(_17341__29_) );
	INVX1 INVX1_2912 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_30_), .Y(_19964_) );
	OAI21X1 OAI21X1_4308 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf0), .B(_19904__bF_buf3), .C(_19153__bF_buf54), .Y(_19965_) );
	AOI21X1 AOI21X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_19964_), .B(_19904__bF_buf2), .C(_19965_), .Y(_17341__30_) );
	INVX1 INVX1_2913 ( .gnd(gnd), .vdd(vdd), .A(registers_a2_31_), .Y(_19966_) );
	OAI21X1 OAI21X1_4309 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf0), .B(_19904__bF_buf1), .C(_19153__bF_buf53), .Y(_19967_) );
	AOI21X1 AOI21X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_19966_), .B(_19904__bF_buf0), .C(_19967_), .Y(_17341__31_) );
	NAND2X1 NAND2X1_3563 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19327_), .Y(_19968_) );
	OAI21X1 OAI21X1_4310 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf52), .Y(_19969_) );
	AOI21X1 AOI21X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_17387_), .B(_19968__bF_buf6), .C(_19969_), .Y(_17340__0_) );
	OAI21X1 OAI21X1_4311 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf51), .Y(_19970_) );
	AOI21X1 AOI21X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_17479_), .B(_19968__bF_buf4), .C(_19970_), .Y(_17340__1_) );
	OAI21X1 OAI21X1_4312 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf50), .Y(_19971_) );
	AOI21X1 AOI21X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_17533_), .B(_19968__bF_buf2), .C(_19971_), .Y(_17340__2_) );
	OAI21X1 OAI21X1_4313 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf49), .Y(_19972_) );
	AOI21X1 AOI21X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_17587_), .B(_19968__bF_buf0), .C(_19972_), .Y(_17340__3_) );
	OAI21X1 OAI21X1_4314 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf48), .Y(_19973_) );
	AOI21X1 AOI21X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_17641_), .B(_19968__bF_buf6), .C(_19973_), .Y(_17340__4_) );
	OAI21X1 OAI21X1_4315 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf47), .Y(_19974_) );
	AOI21X1 AOI21X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_17695_), .B(_19968__bF_buf4), .C(_19974_), .Y(_17340__5_) );
	OAI21X1 OAI21X1_4316 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf46), .Y(_19975_) );
	AOI21X1 AOI21X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_17749_), .B(_19968__bF_buf2), .C(_19975_), .Y(_17340__6_) );
	OAI21X1 OAI21X1_4317 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf45), .Y(_19976_) );
	AOI21X1 AOI21X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_17803_), .B(_19968__bF_buf0), .C(_19976_), .Y(_17340__7_) );
	OAI21X1 OAI21X1_4318 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf44), .Y(_19977_) );
	AOI21X1 AOI21X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_17857_), .B(_19968__bF_buf6), .C(_19977_), .Y(_17340__8_) );
	OAI21X1 OAI21X1_4319 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf43), .Y(_19978_) );
	AOI21X1 AOI21X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_17911_), .B(_19968__bF_buf4), .C(_19978_), .Y(_17340__9_) );
	OAI21X1 OAI21X1_4320 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf42), .Y(_19979_) );
	AOI21X1 AOI21X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_17965_), .B(_19968__bF_buf2), .C(_19979_), .Y(_17340__10_) );
	OAI21X1 OAI21X1_4321 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf41), .Y(_19980_) );
	AOI21X1 AOI21X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_18019_), .B(_19968__bF_buf0), .C(_19980_), .Y(_17340__11_) );
	OAI21X1 OAI21X1_4322 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf40), .Y(_19981_) );
	AOI21X1 AOI21X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_18073_), .B(_19968__bF_buf6), .C(_19981_), .Y(_17340__12_) );
	OAI21X1 OAI21X1_4323 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf39), .Y(_19982_) );
	AOI21X1 AOI21X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_18127_), .B(_19968__bF_buf4), .C(_19982_), .Y(_17340__13_) );
	OAI21X1 OAI21X1_4324 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf38), .Y(_19983_) );
	AOI21X1 AOI21X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_18181_), .B(_19968__bF_buf2), .C(_19983_), .Y(_17340__14_) );
	OAI21X1 OAI21X1_4325 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf37), .Y(_19984_) );
	AOI21X1 AOI21X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_18235_), .B(_19968__bF_buf0), .C(_19984_), .Y(_17340__15_) );
	OAI21X1 OAI21X1_4326 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf36), .Y(_19985_) );
	AOI21X1 AOI21X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_18289_), .B(_19968__bF_buf6), .C(_19985_), .Y(_17340__16_) );
	OAI21X1 OAI21X1_4327 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf35), .Y(_19986_) );
	AOI21X1 AOI21X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_18343_), .B(_19968__bF_buf4), .C(_19986_), .Y(_17340__17_) );
	OAI21X1 OAI21X1_4328 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf34), .Y(_19987_) );
	AOI21X1 AOI21X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_18397_), .B(_19968__bF_buf2), .C(_19987_), .Y(_17340__18_) );
	OAI21X1 OAI21X1_4329 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf33), .Y(_19988_) );
	AOI21X1 AOI21X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_18451_), .B(_19968__bF_buf0), .C(_19988_), .Y(_17340__19_) );
	OAI21X1 OAI21X1_4330 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf32), .Y(_19989_) );
	AOI21X1 AOI21X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_18505_), .B(_19968__bF_buf6), .C(_19989_), .Y(_17340__20_) );
	OAI21X1 OAI21X1_4331 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf31), .Y(_19990_) );
	AOI21X1 AOI21X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_18559_), .B(_19968__bF_buf4), .C(_19990_), .Y(_17340__21_) );
	OAI21X1 OAI21X1_4332 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf30), .Y(_19991_) );
	AOI21X1 AOI21X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_18613_), .B(_19968__bF_buf2), .C(_19991_), .Y(_17340__22_) );
	OAI21X1 OAI21X1_4333 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf29), .Y(_19992_) );
	AOI21X1 AOI21X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_18667_), .B(_19968__bF_buf0), .C(_19992_), .Y(_17340__23_) );
	OAI21X1 OAI21X1_4334 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf28), .Y(_19993_) );
	AOI21X1 AOI21X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_18721_), .B(_19968__bF_buf6), .C(_19993_), .Y(_17340__24_) );
	OAI21X1 OAI21X1_4335 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf27), .Y(_19994_) );
	AOI21X1 AOI21X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_18775_), .B(_19968__bF_buf4), .C(_19994_), .Y(_17340__25_) );
	OAI21X1 OAI21X1_4336 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf26), .Y(_19995_) );
	AOI21X1 AOI21X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_18829_), .B(_19968__bF_buf2), .C(_19995_), .Y(_17340__26_) );
	OAI21X1 OAI21X1_4337 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf25), .Y(_19996_) );
	AOI21X1 AOI21X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_18883_), .B(_19968__bF_buf0), .C(_19996_), .Y(_17340__27_) );
	OAI21X1 OAI21X1_4338 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_19968__bF_buf7), .C(_19153__bF_buf24), .Y(_19997_) );
	AOI21X1 AOI21X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_18937_), .B(_19968__bF_buf6), .C(_19997_), .Y(_17340__28_) );
	OAI21X1 OAI21X1_4339 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_19968__bF_buf5), .C(_19153__bF_buf23), .Y(_19998_) );
	AOI21X1 AOI21X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_18991_), .B(_19968__bF_buf4), .C(_19998_), .Y(_17340__29_) );
	OAI21X1 OAI21X1_4340 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_19968__bF_buf3), .C(_19153__bF_buf22), .Y(_19999_) );
	AOI21X1 AOI21X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_19045_), .B(_19968__bF_buf2), .C(_19999_), .Y(_17340__30_) );
	OAI21X1 OAI21X1_4341 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_19968__bF_buf1), .C(_19153__bF_buf21), .Y(_20000_) );
	AOI21X1 AOI21X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_19099_), .B(_19968__bF_buf0), .C(_20000_), .Y(_17340__31_) );
	INVX1 INVX1_2914 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_0_), .Y(_20001_) );
	NAND2X1 NAND2X1_3564 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19361_), .Y(_20002_) );
	OAI21X1 OAI21X1_4342 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf20), .Y(_20003_) );
	AOI21X1 AOI21X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_20001_), .B(_20002__bF_buf6), .C(_20003_), .Y(_17339__0_) );
	INVX1 INVX1_2915 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_1_), .Y(_20004_) );
	OAI21X1 OAI21X1_4343 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf19), .Y(_20005_) );
	AOI21X1 AOI21X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_20004_), .B(_20002__bF_buf4), .C(_20005_), .Y(_17339__1_) );
	INVX1 INVX1_2916 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_2_), .Y(_20006_) );
	OAI21X1 OAI21X1_4344 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf18), .Y(_20007_) );
	AOI21X1 AOI21X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_20006_), .B(_20002__bF_buf2), .C(_20007_), .Y(_17339__2_) );
	INVX1 INVX1_2917 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_3_), .Y(_20008_) );
	OAI21X1 OAI21X1_4345 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf17), .Y(_20009_) );
	AOI21X1 AOI21X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_20008_), .B(_20002__bF_buf0), .C(_20009_), .Y(_17339__3_) );
	INVX1 INVX1_2918 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_4_), .Y(_20010_) );
	OAI21X1 OAI21X1_4346 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf16), .Y(_20011_) );
	AOI21X1 AOI21X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_20010_), .B(_20002__bF_buf6), .C(_20011_), .Y(_17339__4_) );
	INVX1 INVX1_2919 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_5_), .Y(_20012_) );
	OAI21X1 OAI21X1_4347 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf15), .Y(_20013_) );
	AOI21X1 AOI21X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_20012_), .B(_20002__bF_buf4), .C(_20013_), .Y(_17339__5_) );
	INVX1 INVX1_2920 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_6_), .Y(_20014_) );
	OAI21X1 OAI21X1_4348 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf14), .Y(_20015_) );
	AOI21X1 AOI21X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_20014_), .B(_20002__bF_buf2), .C(_20015_), .Y(_17339__6_) );
	INVX1 INVX1_2921 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_7_), .Y(_20016_) );
	OAI21X1 OAI21X1_4349 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf13), .Y(_20017_) );
	AOI21X1 AOI21X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_20016_), .B(_20002__bF_buf0), .C(_20017_), .Y(_17339__7_) );
	INVX1 INVX1_2922 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_8_), .Y(_20018_) );
	OAI21X1 OAI21X1_4350 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf12), .Y(_20019_) );
	AOI21X1 AOI21X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_20018_), .B(_20002__bF_buf6), .C(_20019_), .Y(_17339__8_) );
	INVX1 INVX1_2923 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_9_), .Y(_20020_) );
	OAI21X1 OAI21X1_4351 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf11), .Y(_20021_) );
	AOI21X1 AOI21X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_20020_), .B(_20002__bF_buf4), .C(_20021_), .Y(_17339__9_) );
	INVX1 INVX1_2924 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_10_), .Y(_20022_) );
	OAI21X1 OAI21X1_4352 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf10), .Y(_20023_) );
	AOI21X1 AOI21X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_20022_), .B(_20002__bF_buf2), .C(_20023_), .Y(_17339__10_) );
	INVX1 INVX1_2925 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_11_), .Y(_20024_) );
	OAI21X1 OAI21X1_4353 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf9), .Y(_20025_) );
	AOI21X1 AOI21X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_20024_), .B(_20002__bF_buf0), .C(_20025_), .Y(_17339__11_) );
	INVX1 INVX1_2926 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_12_), .Y(_20026_) );
	OAI21X1 OAI21X1_4354 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf8), .Y(_20027_) );
	AOI21X1 AOI21X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_20026_), .B(_20002__bF_buf6), .C(_20027_), .Y(_17339__12_) );
	INVX1 INVX1_2927 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_13_), .Y(_20028_) );
	OAI21X1 OAI21X1_4355 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf7), .Y(_20029_) );
	AOI21X1 AOI21X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_20028_), .B(_20002__bF_buf4), .C(_20029_), .Y(_17339__13_) );
	INVX1 INVX1_2928 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_14_), .Y(_20030_) );
	OAI21X1 OAI21X1_4356 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf6), .Y(_20031_) );
	AOI21X1 AOI21X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_20030_), .B(_20002__bF_buf2), .C(_20031_), .Y(_17339__14_) );
	INVX1 INVX1_2929 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_15_), .Y(_20032_) );
	OAI21X1 OAI21X1_4357 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf5), .Y(_20033_) );
	AOI21X1 AOI21X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_20032_), .B(_20002__bF_buf0), .C(_20033_), .Y(_17339__15_) );
	INVX1 INVX1_2930 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_16_), .Y(_20034_) );
	OAI21X1 OAI21X1_4358 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf4), .Y(_20035_) );
	AOI21X1 AOI21X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_20034_), .B(_20002__bF_buf6), .C(_20035_), .Y(_17339__16_) );
	INVX1 INVX1_2931 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_17_), .Y(_20036_) );
	OAI21X1 OAI21X1_4359 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf3), .Y(_20037_) );
	AOI21X1 AOI21X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_20036_), .B(_20002__bF_buf4), .C(_20037_), .Y(_17339__17_) );
	INVX1 INVX1_2932 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_18_), .Y(_20038_) );
	OAI21X1 OAI21X1_4360 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf2), .Y(_20039_) );
	AOI21X1 AOI21X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_20038_), .B(_20002__bF_buf2), .C(_20039_), .Y(_17339__18_) );
	INVX1 INVX1_2933 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_19_), .Y(_20040_) );
	OAI21X1 OAI21X1_4361 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf1), .Y(_20041_) );
	AOI21X1 AOI21X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_20040_), .B(_20002__bF_buf0), .C(_20041_), .Y(_17339__19_) );
	INVX1 INVX1_2934 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_20_), .Y(_20042_) );
	OAI21X1 OAI21X1_4362 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf0), .Y(_20043_) );
	AOI21X1 AOI21X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_20042_), .B(_20002__bF_buf6), .C(_20043_), .Y(_17339__20_) );
	INVX1 INVX1_2935 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_21_), .Y(_20044_) );
	OAI21X1 OAI21X1_4363 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf98), .Y(_20045_) );
	AOI21X1 AOI21X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_20044_), .B(_20002__bF_buf4), .C(_20045_), .Y(_17339__21_) );
	INVX1 INVX1_2936 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_22_), .Y(_20046_) );
	OAI21X1 OAI21X1_4364 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf97), .Y(_20047_) );
	AOI21X1 AOI21X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_20046_), .B(_20002__bF_buf2), .C(_20047_), .Y(_17339__22_) );
	INVX1 INVX1_2937 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_23_), .Y(_20048_) );
	OAI21X1 OAI21X1_4365 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf96), .Y(_20049_) );
	AOI21X1 AOI21X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_20048_), .B(_20002__bF_buf0), .C(_20049_), .Y(_17339__23_) );
	INVX1 INVX1_2938 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_24_), .Y(_20050_) );
	OAI21X1 OAI21X1_4366 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf95), .Y(_20051_) );
	AOI21X1 AOI21X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_20050_), .B(_20002__bF_buf6), .C(_20051_), .Y(_17339__24_) );
	INVX1 INVX1_2939 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_25_), .Y(_20052_) );
	OAI21X1 OAI21X1_4367 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf94), .Y(_20053_) );
	AOI21X1 AOI21X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_20052_), .B(_20002__bF_buf4), .C(_20053_), .Y(_17339__25_) );
	INVX1 INVX1_2940 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_26_), .Y(_20054_) );
	OAI21X1 OAI21X1_4368 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf93), .Y(_20055_) );
	AOI21X1 AOI21X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_20054_), .B(_20002__bF_buf2), .C(_20055_), .Y(_17339__26_) );
	INVX1 INVX1_2941 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_27_), .Y(_20056_) );
	OAI21X1 OAI21X1_4369 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf92), .Y(_20057_) );
	AOI21X1 AOI21X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_20056_), .B(_20002__bF_buf0), .C(_20057_), .Y(_17339__27_) );
	INVX1 INVX1_2942 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_28_), .Y(_20058_) );
	OAI21X1 OAI21X1_4370 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf3), .B(_20002__bF_buf7), .C(_19153__bF_buf91), .Y(_20059_) );
	AOI21X1 AOI21X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_20058_), .B(_20002__bF_buf6), .C(_20059_), .Y(_17339__28_) );
	INVX1 INVX1_2943 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_29_), .Y(_20060_) );
	OAI21X1 OAI21X1_4371 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf3), .B(_20002__bF_buf5), .C(_19153__bF_buf90), .Y(_20061_) );
	AOI21X1 AOI21X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_20060_), .B(_20002__bF_buf4), .C(_20061_), .Y(_17339__29_) );
	INVX1 INVX1_2944 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_30_), .Y(_20062_) );
	OAI21X1 OAI21X1_4372 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf3), .B(_20002__bF_buf3), .C(_19153__bF_buf89), .Y(_20063_) );
	AOI21X1 AOI21X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_20062_), .B(_20002__bF_buf2), .C(_20063_), .Y(_17339__30_) );
	INVX1 INVX1_2945 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_31_), .Y(_20064_) );
	OAI21X1 OAI21X1_4373 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf3), .B(_20002__bF_buf1), .C(_19153__bF_buf88), .Y(_20065_) );
	AOI21X1 AOI21X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_20064_), .B(_20002__bF_buf0), .C(_20065_), .Y(_17339__31_) );
	NAND2X1 NAND2X1_3565 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19395_), .Y(_20066_) );
	OAI21X1 OAI21X1_4374 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf87), .Y(_20067_) );
	AOI21X1 AOI21X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_17388_), .B(_20066__bF_buf6), .C(_20067_), .Y(_17369__0_) );
	OAI21X1 OAI21X1_4375 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf86), .Y(_20068_) );
	AOI21X1 AOI21X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_17480_), .B(_20066__bF_buf4), .C(_20068_), .Y(_17369__1_) );
	OAI21X1 OAI21X1_4376 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf85), .Y(_20069_) );
	AOI21X1 AOI21X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_17534_), .B(_20066__bF_buf2), .C(_20069_), .Y(_17369__2_) );
	OAI21X1 OAI21X1_4377 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf84), .Y(_20070_) );
	AOI21X1 AOI21X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_17588_), .B(_20066__bF_buf0), .C(_20070_), .Y(_17369__3_) );
	OAI21X1 OAI21X1_4378 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf83), .Y(_20071_) );
	AOI21X1 AOI21X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_17642_), .B(_20066__bF_buf6), .C(_20071_), .Y(_17369__4_) );
	OAI21X1 OAI21X1_4379 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf82), .Y(_20072_) );
	AOI21X1 AOI21X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_17696_), .B(_20066__bF_buf4), .C(_20072_), .Y(_17369__5_) );
	OAI21X1 OAI21X1_4380 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf81), .Y(_20073_) );
	AOI21X1 AOI21X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_17750_), .B(_20066__bF_buf2), .C(_20073_), .Y(_17369__6_) );
	OAI21X1 OAI21X1_4381 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf80), .Y(_20074_) );
	AOI21X1 AOI21X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_17804_), .B(_20066__bF_buf0), .C(_20074_), .Y(_17369__7_) );
	OAI21X1 OAI21X1_4382 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf79), .Y(_20075_) );
	AOI21X1 AOI21X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_17858_), .B(_20066__bF_buf6), .C(_20075_), .Y(_17369__8_) );
	OAI21X1 OAI21X1_4383 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf78), .Y(_20076_) );
	AOI21X1 AOI21X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_17912_), .B(_20066__bF_buf4), .C(_20076_), .Y(_17369__9_) );
	OAI21X1 OAI21X1_4384 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf77), .Y(_20077_) );
	AOI21X1 AOI21X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_17966_), .B(_20066__bF_buf2), .C(_20077_), .Y(_17369__10_) );
	OAI21X1 OAI21X1_4385 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf76), .Y(_20078_) );
	AOI21X1 AOI21X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_18020_), .B(_20066__bF_buf0), .C(_20078_), .Y(_17369__11_) );
	OAI21X1 OAI21X1_4386 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf75), .Y(_20079_) );
	AOI21X1 AOI21X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_18074_), .B(_20066__bF_buf6), .C(_20079_), .Y(_17369__12_) );
	OAI21X1 OAI21X1_4387 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf74), .Y(_20080_) );
	AOI21X1 AOI21X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_18128_), .B(_20066__bF_buf4), .C(_20080_), .Y(_17369__13_) );
	OAI21X1 OAI21X1_4388 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf73), .Y(_20081_) );
	AOI21X1 AOI21X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_18182_), .B(_20066__bF_buf2), .C(_20081_), .Y(_17369__14_) );
	OAI21X1 OAI21X1_4389 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf72), .Y(_20082_) );
	AOI21X1 AOI21X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_18236_), .B(_20066__bF_buf0), .C(_20082_), .Y(_17369__15_) );
	OAI21X1 OAI21X1_4390 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf71), .Y(_20083_) );
	AOI21X1 AOI21X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_18290_), .B(_20066__bF_buf6), .C(_20083_), .Y(_17369__16_) );
	OAI21X1 OAI21X1_4391 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf70), .Y(_20084_) );
	AOI21X1 AOI21X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_18344_), .B(_20066__bF_buf4), .C(_20084_), .Y(_17369__17_) );
	OAI21X1 OAI21X1_4392 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf69), .Y(_20085_) );
	AOI21X1 AOI21X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_18398_), .B(_20066__bF_buf2), .C(_20085_), .Y(_17369__18_) );
	OAI21X1 OAI21X1_4393 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf68), .Y(_20086_) );
	AOI21X1 AOI21X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_18452_), .B(_20066__bF_buf0), .C(_20086_), .Y(_17369__19_) );
	OAI21X1 OAI21X1_4394 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf67), .Y(_20087_) );
	AOI21X1 AOI21X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_18506_), .B(_20066__bF_buf6), .C(_20087_), .Y(_17369__20_) );
	OAI21X1 OAI21X1_4395 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf66), .Y(_20088_) );
	AOI21X1 AOI21X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_18560_), .B(_20066__bF_buf4), .C(_20088_), .Y(_17369__21_) );
	OAI21X1 OAI21X1_4396 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf65), .Y(_20089_) );
	AOI21X1 AOI21X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_18614_), .B(_20066__bF_buf2), .C(_20089_), .Y(_17369__22_) );
	OAI21X1 OAI21X1_4397 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf64), .Y(_20090_) );
	AOI21X1 AOI21X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_18668_), .B(_20066__bF_buf0), .C(_20090_), .Y(_17369__23_) );
	OAI21X1 OAI21X1_4398 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf63), .Y(_20091_) );
	AOI21X1 AOI21X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_18722_), .B(_20066__bF_buf6), .C(_20091_), .Y(_17369__24_) );
	OAI21X1 OAI21X1_4399 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf62), .Y(_20092_) );
	AOI21X1 AOI21X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_18776_), .B(_20066__bF_buf4), .C(_20092_), .Y(_17369__25_) );
	OAI21X1 OAI21X1_4400 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf61), .Y(_20093_) );
	AOI21X1 AOI21X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_18830_), .B(_20066__bF_buf2), .C(_20093_), .Y(_17369__26_) );
	OAI21X1 OAI21X1_4401 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf60), .Y(_20094_) );
	AOI21X1 AOI21X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_18884_), .B(_20066__bF_buf0), .C(_20094_), .Y(_17369__27_) );
	OAI21X1 OAI21X1_4402 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf2), .B(_20066__bF_buf7), .C(_19153__bF_buf59), .Y(_20095_) );
	AOI21X1 AOI21X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_18938_), .B(_20066__bF_buf6), .C(_20095_), .Y(_17369__28_) );
	OAI21X1 OAI21X1_4403 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf2), .B(_20066__bF_buf5), .C(_19153__bF_buf58), .Y(_20096_) );
	AOI21X1 AOI21X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_18992_), .B(_20066__bF_buf4), .C(_20096_), .Y(_17369__29_) );
	OAI21X1 OAI21X1_4404 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf2), .B(_20066__bF_buf3), .C(_19153__bF_buf57), .Y(_20097_) );
	AOI21X1 AOI21X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_19046_), .B(_20066__bF_buf2), .C(_20097_), .Y(_17369__30_) );
	OAI21X1 OAI21X1_4405 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf2), .B(_20066__bF_buf1), .C(_19153__bF_buf56), .Y(_20098_) );
	AOI21X1 AOI21X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_19100_), .B(_20066__bF_buf0), .C(_20098_), .Y(_17369__31_) );
	INVX1 INVX1_2946 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_0_), .Y(_20099_) );
	AND2X2 AND2X2_421 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19289_), .Y(_20100_) );
	NAND2X1 NAND2X1_3566 ( .gnd(gnd), .vdd(vdd), .A(_19431_), .B(_20100_), .Y(_20101_) );
	OAI21X1 OAI21X1_4406 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf55), .Y(_20102_) );
	AOI21X1 AOI21X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_20099_), .B(_20101__bF_buf6), .C(_20102_), .Y(_17368__0_) );
	INVX1 INVX1_2947 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_1_), .Y(_20103_) );
	OAI21X1 OAI21X1_4407 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf54), .Y(_20104_) );
	AOI21X1 AOI21X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_20103_), .B(_20101__bF_buf4), .C(_20104_), .Y(_17368__1_) );
	INVX1 INVX1_2948 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_2_), .Y(_20105_) );
	OAI21X1 OAI21X1_4408 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf53), .Y(_20106_) );
	AOI21X1 AOI21X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_20105_), .B(_20101__bF_buf2), .C(_20106_), .Y(_17368__2_) );
	INVX1 INVX1_2949 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_3_), .Y(_20107_) );
	OAI21X1 OAI21X1_4409 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf52), .Y(_20108_) );
	AOI21X1 AOI21X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_20107_), .B(_20101__bF_buf0), .C(_20108_), .Y(_17368__3_) );
	INVX1 INVX1_2950 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_4_), .Y(_20109_) );
	OAI21X1 OAI21X1_4410 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf51), .Y(_20110_) );
	AOI21X1 AOI21X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_20109_), .B(_20101__bF_buf6), .C(_20110_), .Y(_17368__4_) );
	INVX1 INVX1_2951 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_5_), .Y(_20111_) );
	OAI21X1 OAI21X1_4411 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf50), .Y(_20112_) );
	AOI21X1 AOI21X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_20111_), .B(_20101__bF_buf4), .C(_20112_), .Y(_17368__5_) );
	INVX1 INVX1_2952 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_6_), .Y(_20113_) );
	OAI21X1 OAI21X1_4412 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf49), .Y(_20114_) );
	AOI21X1 AOI21X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_20113_), .B(_20101__bF_buf2), .C(_20114_), .Y(_17368__6_) );
	INVX1 INVX1_2953 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_7_), .Y(_20115_) );
	OAI21X1 OAI21X1_4413 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf48), .Y(_20116_) );
	AOI21X1 AOI21X1_2898 ( .gnd(gnd), .vdd(vdd), .A(_20115_), .B(_20101__bF_buf0), .C(_20116_), .Y(_17368__7_) );
	INVX1 INVX1_2954 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_8_), .Y(_20117_) );
	OAI21X1 OAI21X1_4414 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf47), .Y(_20118_) );
	AOI21X1 AOI21X1_2899 ( .gnd(gnd), .vdd(vdd), .A(_20117_), .B(_20101__bF_buf6), .C(_20118_), .Y(_17368__8_) );
	INVX1 INVX1_2955 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_9_), .Y(_20119_) );
	OAI21X1 OAI21X1_4415 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf46), .Y(_20120_) );
	AOI21X1 AOI21X1_2900 ( .gnd(gnd), .vdd(vdd), .A(_20119_), .B(_20101__bF_buf4), .C(_20120_), .Y(_17368__9_) );
	INVX1 INVX1_2956 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_10_), .Y(_20121_) );
	OAI21X1 OAI21X1_4416 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf45), .Y(_20122_) );
	AOI21X1 AOI21X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_20121_), .B(_20101__bF_buf2), .C(_20122_), .Y(_17368__10_) );
	INVX1 INVX1_2957 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_11_), .Y(_20123_) );
	OAI21X1 OAI21X1_4417 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf44), .Y(_20124_) );
	AOI21X1 AOI21X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_20123_), .B(_20101__bF_buf0), .C(_20124_), .Y(_17368__11_) );
	INVX1 INVX1_2958 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_12_), .Y(_20125_) );
	OAI21X1 OAI21X1_4418 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf43), .Y(_20126_) );
	AOI21X1 AOI21X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_20125_), .B(_20101__bF_buf6), .C(_20126_), .Y(_17368__12_) );
	INVX1 INVX1_2959 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_13_), .Y(_20127_) );
	OAI21X1 OAI21X1_4419 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf42), .Y(_20128_) );
	AOI21X1 AOI21X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_20127_), .B(_20101__bF_buf4), .C(_20128_), .Y(_17368__13_) );
	INVX1 INVX1_2960 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_14_), .Y(_20129_) );
	OAI21X1 OAI21X1_4420 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf41), .Y(_20130_) );
	AOI21X1 AOI21X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_20129_), .B(_20101__bF_buf2), .C(_20130_), .Y(_17368__14_) );
	INVX1 INVX1_2961 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_15_), .Y(_20131_) );
	OAI21X1 OAI21X1_4421 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf40), .Y(_20132_) );
	AOI21X1 AOI21X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_20131_), .B(_20101__bF_buf0), .C(_20132_), .Y(_17368__15_) );
	INVX1 INVX1_2962 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_16_), .Y(_20133_) );
	OAI21X1 OAI21X1_4422 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf39), .Y(_20134_) );
	AOI21X1 AOI21X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_20133_), .B(_20101__bF_buf6), .C(_20134_), .Y(_17368__16_) );
	INVX1 INVX1_2963 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_17_), .Y(_20135_) );
	OAI21X1 OAI21X1_4423 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf38), .Y(_20136_) );
	AOI21X1 AOI21X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_20135_), .B(_20101__bF_buf4), .C(_20136_), .Y(_17368__17_) );
	INVX1 INVX1_2964 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_18_), .Y(_20137_) );
	OAI21X1 OAI21X1_4424 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf37), .Y(_20138_) );
	AOI21X1 AOI21X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_20137_), .B(_20101__bF_buf2), .C(_20138_), .Y(_17368__18_) );
	INVX1 INVX1_2965 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_19_), .Y(_20139_) );
	OAI21X1 OAI21X1_4425 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf36), .Y(_20140_) );
	AOI21X1 AOI21X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_20139_), .B(_20101__bF_buf0), .C(_20140_), .Y(_17368__19_) );
	INVX1 INVX1_2966 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_20_), .Y(_20141_) );
	OAI21X1 OAI21X1_4426 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf35), .Y(_20142_) );
	AOI21X1 AOI21X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_20141_), .B(_20101__bF_buf6), .C(_20142_), .Y(_17368__20_) );
	INVX1 INVX1_2967 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_21_), .Y(_20143_) );
	OAI21X1 OAI21X1_4427 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf34), .Y(_20144_) );
	AOI21X1 AOI21X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_20143_), .B(_20101__bF_buf4), .C(_20144_), .Y(_17368__21_) );
	INVX1 INVX1_2968 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_22_), .Y(_20145_) );
	OAI21X1 OAI21X1_4428 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf33), .Y(_20146_) );
	AOI21X1 AOI21X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_20145_), .B(_20101__bF_buf2), .C(_20146_), .Y(_17368__22_) );
	INVX1 INVX1_2969 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_23_), .Y(_20147_) );
	OAI21X1 OAI21X1_4429 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf32), .Y(_20148_) );
	AOI21X1 AOI21X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_20147_), .B(_20101__bF_buf0), .C(_20148_), .Y(_17368__23_) );
	INVX1 INVX1_2970 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_24_), .Y(_20149_) );
	OAI21X1 OAI21X1_4430 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf31), .Y(_20150_) );
	AOI21X1 AOI21X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_20149_), .B(_20101__bF_buf6), .C(_20150_), .Y(_17368__24_) );
	INVX1 INVX1_2971 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_25_), .Y(_20151_) );
	OAI21X1 OAI21X1_4431 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf30), .Y(_20152_) );
	AOI21X1 AOI21X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_20151_), .B(_20101__bF_buf4), .C(_20152_), .Y(_17368__25_) );
	INVX1 INVX1_2972 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_26_), .Y(_20153_) );
	OAI21X1 OAI21X1_4432 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf29), .Y(_20154_) );
	AOI21X1 AOI21X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_20153_), .B(_20101__bF_buf2), .C(_20154_), .Y(_17368__26_) );
	INVX1 INVX1_2973 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_27_), .Y(_20155_) );
	OAI21X1 OAI21X1_4433 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf28), .Y(_20156_) );
	AOI21X1 AOI21X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_20155_), .B(_20101__bF_buf0), .C(_20156_), .Y(_17368__27_) );
	INVX1 INVX1_2974 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_28_), .Y(_20157_) );
	OAI21X1 OAI21X1_4434 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf1), .B(_20101__bF_buf7), .C(_19153__bF_buf27), .Y(_20158_) );
	AOI21X1 AOI21X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_20157_), .B(_20101__bF_buf6), .C(_20158_), .Y(_17368__28_) );
	INVX1 INVX1_2975 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_29_), .Y(_20159_) );
	OAI21X1 OAI21X1_4435 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf1), .B(_20101__bF_buf5), .C(_19153__bF_buf26), .Y(_20160_) );
	AOI21X1 AOI21X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_20159_), .B(_20101__bF_buf4), .C(_20160_), .Y(_17368__29_) );
	INVX1 INVX1_2976 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_30_), .Y(_20161_) );
	OAI21X1 OAI21X1_4436 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf1), .B(_20101__bF_buf3), .C(_19153__bF_buf25), .Y(_20162_) );
	AOI21X1 AOI21X1_2921 ( .gnd(gnd), .vdd(vdd), .A(_20161_), .B(_20101__bF_buf2), .C(_20162_), .Y(_17368__30_) );
	INVX1 INVX1_2977 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_31_), .Y(_20163_) );
	OAI21X1 OAI21X1_4437 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf1), .B(_20101__bF_buf1), .C(_19153__bF_buf24), .Y(_20164_) );
	AOI21X1 AOI21X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_20163_), .B(_20101__bF_buf0), .C(_20164_), .Y(_17368__31_) );
	INVX1 INVX1_2978 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_0_), .Y(_20165_) );
	NAND2X1 NAND2X1_3567 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19498_), .Y(_20166_) );
	OAI21X1 OAI21X1_4438 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf23), .Y(_20167_) );
	AOI21X1 AOI21X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_20165_), .B(_20166__bF_buf6), .C(_20167_), .Y(_17367__0_) );
	INVX1 INVX1_2979 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_1_), .Y(_20168_) );
	OAI21X1 OAI21X1_4439 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf22), .Y(_20169_) );
	AOI21X1 AOI21X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_20168_), .B(_20166__bF_buf4), .C(_20169_), .Y(_17367__1_) );
	INVX1 INVX1_2980 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_2_), .Y(_20170_) );
	OAI21X1 OAI21X1_4440 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf21), .Y(_20171_) );
	AOI21X1 AOI21X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_20170_), .B(_20166__bF_buf2), .C(_20171_), .Y(_17367__2_) );
	INVX1 INVX1_2981 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_3_), .Y(_20172_) );
	OAI21X1 OAI21X1_4441 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf20), .Y(_20173_) );
	AOI21X1 AOI21X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_20172_), .B(_20166__bF_buf0), .C(_20173_), .Y(_17367__3_) );
	INVX1 INVX1_2982 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_4_), .Y(_20174_) );
	OAI21X1 OAI21X1_4442 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf19), .Y(_20175_) );
	AOI21X1 AOI21X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_20174_), .B(_20166__bF_buf6), .C(_20175_), .Y(_17367__4_) );
	INVX1 INVX1_2983 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_5_), .Y(_20176_) );
	OAI21X1 OAI21X1_4443 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf18), .Y(_20177_) );
	AOI21X1 AOI21X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_20176_), .B(_20166__bF_buf4), .C(_20177_), .Y(_17367__5_) );
	INVX1 INVX1_2984 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_6_), .Y(_20178_) );
	OAI21X1 OAI21X1_4444 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf17), .Y(_20179_) );
	AOI21X1 AOI21X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_20178_), .B(_20166__bF_buf2), .C(_20179_), .Y(_17367__6_) );
	INVX1 INVX1_2985 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_7_), .Y(_20180_) );
	OAI21X1 OAI21X1_4445 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf16), .Y(_20181_) );
	AOI21X1 AOI21X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_20180_), .B(_20166__bF_buf0), .C(_20181_), .Y(_17367__7_) );
	INVX1 INVX1_2986 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_8_), .Y(_20182_) );
	OAI21X1 OAI21X1_4446 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf15), .Y(_20183_) );
	AOI21X1 AOI21X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_20182_), .B(_20166__bF_buf6), .C(_20183_), .Y(_17367__8_) );
	INVX1 INVX1_2987 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_9_), .Y(_20184_) );
	OAI21X1 OAI21X1_4447 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf14), .Y(_20185_) );
	AOI21X1 AOI21X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_20184_), .B(_20166__bF_buf4), .C(_20185_), .Y(_17367__9_) );
	INVX1 INVX1_2988 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_10_), .Y(_20186_) );
	OAI21X1 OAI21X1_4448 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf13), .Y(_20187_) );
	AOI21X1 AOI21X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_20186_), .B(_20166__bF_buf2), .C(_20187_), .Y(_17367__10_) );
	INVX1 INVX1_2989 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_11_), .Y(_20188_) );
	OAI21X1 OAI21X1_4449 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf12), .Y(_20189_) );
	AOI21X1 AOI21X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_20188_), .B(_20166__bF_buf0), .C(_20189_), .Y(_17367__11_) );
	INVX1 INVX1_2990 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_12_), .Y(_20190_) );
	OAI21X1 OAI21X1_4450 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf11), .Y(_20191_) );
	AOI21X1 AOI21X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_20190_), .B(_20166__bF_buf6), .C(_20191_), .Y(_17367__12_) );
	INVX1 INVX1_2991 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_13_), .Y(_20192_) );
	OAI21X1 OAI21X1_4451 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf10), .Y(_20193_) );
	AOI21X1 AOI21X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_20192_), .B(_20166__bF_buf4), .C(_20193_), .Y(_17367__13_) );
	INVX1 INVX1_2992 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_14_), .Y(_20194_) );
	OAI21X1 OAI21X1_4452 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf9), .Y(_20195_) );
	AOI21X1 AOI21X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_20194_), .B(_20166__bF_buf2), .C(_20195_), .Y(_17367__14_) );
	INVX1 INVX1_2993 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_15_), .Y(_20196_) );
	OAI21X1 OAI21X1_4453 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf8), .Y(_20197_) );
	AOI21X1 AOI21X1_2938 ( .gnd(gnd), .vdd(vdd), .A(_20196_), .B(_20166__bF_buf0), .C(_20197_), .Y(_17367__15_) );
	INVX1 INVX1_2994 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_16_), .Y(_20198_) );
	OAI21X1 OAI21X1_4454 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf7), .Y(_20199_) );
	AOI21X1 AOI21X1_2939 ( .gnd(gnd), .vdd(vdd), .A(_20198_), .B(_20166__bF_buf6), .C(_20199_), .Y(_17367__16_) );
	INVX1 INVX1_2995 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_17_), .Y(_20200_) );
	OAI21X1 OAI21X1_4455 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf6), .Y(_20201_) );
	AOI21X1 AOI21X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_20200_), .B(_20166__bF_buf4), .C(_20201_), .Y(_17367__17_) );
	INVX1 INVX1_2996 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_18_), .Y(_20202_) );
	OAI21X1 OAI21X1_4456 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf5), .Y(_20203_) );
	AOI21X1 AOI21X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_20202_), .B(_20166__bF_buf2), .C(_20203_), .Y(_17367__18_) );
	INVX1 INVX1_2997 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_19_), .Y(_20204_) );
	OAI21X1 OAI21X1_4457 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf4), .Y(_20205_) );
	AOI21X1 AOI21X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_20204_), .B(_20166__bF_buf0), .C(_20205_), .Y(_17367__19_) );
	INVX1 INVX1_2998 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_20_), .Y(_20206_) );
	OAI21X1 OAI21X1_4458 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf3), .Y(_20207_) );
	AOI21X1 AOI21X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_20206_), .B(_20166__bF_buf6), .C(_20207_), .Y(_17367__20_) );
	INVX1 INVX1_2999 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_21_), .Y(_20208_) );
	OAI21X1 OAI21X1_4459 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf2), .Y(_20209_) );
	AOI21X1 AOI21X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_20208_), .B(_20166__bF_buf4), .C(_20209_), .Y(_17367__21_) );
	INVX1 INVX1_3000 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_22_), .Y(_20210_) );
	OAI21X1 OAI21X1_4460 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf1), .Y(_20211_) );
	AOI21X1 AOI21X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_20210_), .B(_20166__bF_buf2), .C(_20211_), .Y(_17367__22_) );
	INVX1 INVX1_3001 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_23_), .Y(_20212_) );
	OAI21X1 OAI21X1_4461 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf0), .Y(_20213_) );
	AOI21X1 AOI21X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_20212_), .B(_20166__bF_buf0), .C(_20213_), .Y(_17367__23_) );
	INVX1 INVX1_3002 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_24_), .Y(_20214_) );
	OAI21X1 OAI21X1_4462 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf98), .Y(_20215_) );
	AOI21X1 AOI21X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_20214_), .B(_20166__bF_buf6), .C(_20215_), .Y(_17367__24_) );
	INVX1 INVX1_3003 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_25_), .Y(_20216_) );
	OAI21X1 OAI21X1_4463 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf97), .Y(_20217_) );
	AOI21X1 AOI21X1_2948 ( .gnd(gnd), .vdd(vdd), .A(_20216_), .B(_20166__bF_buf4), .C(_20217_), .Y(_17367__25_) );
	INVX1 INVX1_3004 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_26_), .Y(_20218_) );
	OAI21X1 OAI21X1_4464 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf96), .Y(_20219_) );
	AOI21X1 AOI21X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_20218_), .B(_20166__bF_buf2), .C(_20219_), .Y(_17367__26_) );
	INVX1 INVX1_3005 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_27_), .Y(_20220_) );
	OAI21X1 OAI21X1_4465 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf95), .Y(_20221_) );
	AOI21X1 AOI21X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_20220_), .B(_20166__bF_buf0), .C(_20221_), .Y(_17367__27_) );
	INVX1 INVX1_3006 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_28_), .Y(_20222_) );
	OAI21X1 OAI21X1_4466 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf0), .B(_20166__bF_buf7), .C(_19153__bF_buf94), .Y(_20223_) );
	AOI21X1 AOI21X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_20222_), .B(_20166__bF_buf6), .C(_20223_), .Y(_17367__28_) );
	INVX1 INVX1_3007 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_29_), .Y(_20224_) );
	OAI21X1 OAI21X1_4467 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf0), .B(_20166__bF_buf5), .C(_19153__bF_buf93), .Y(_20225_) );
	AOI21X1 AOI21X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_20224_), .B(_20166__bF_buf4), .C(_20225_), .Y(_17367__29_) );
	INVX1 INVX1_3008 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_30_), .Y(_20226_) );
	OAI21X1 OAI21X1_4468 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf0), .B(_20166__bF_buf3), .C(_19153__bF_buf92), .Y(_20227_) );
	AOI21X1 AOI21X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_20226_), .B(_20166__bF_buf2), .C(_20227_), .Y(_17367__30_) );
	INVX1 INVX1_3009 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_31_), .Y(_20228_) );
	OAI21X1 OAI21X1_4469 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf0), .B(_20166__bF_buf1), .C(_19153__bF_buf91), .Y(_20229_) );
	AOI21X1 AOI21X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_20228_), .B(_20166__bF_buf0), .C(_20229_), .Y(_17367__31_) );
	INVX1 INVX1_3010 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_0_), .Y(_20230_) );
	NAND2X1 NAND2X1_3568 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19532_), .Y(_20231_) );
	OAI21X1 OAI21X1_4470 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf90), .Y(_20232_) );
	AOI21X1 AOI21X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_20230_), .B(_20231__bF_buf6), .C(_20232_), .Y(_17366__0_) );
	INVX1 INVX1_3011 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_1_), .Y(_20233_) );
	OAI21X1 OAI21X1_4471 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf89), .Y(_20234_) );
	AOI21X1 AOI21X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_20233_), .B(_20231__bF_buf4), .C(_20234_), .Y(_17366__1_) );
	INVX1 INVX1_3012 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_2_), .Y(_20235_) );
	OAI21X1 OAI21X1_4472 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf88), .Y(_20236_) );
	AOI21X1 AOI21X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_20235_), .B(_20231__bF_buf2), .C(_20236_), .Y(_17366__2_) );
	INVX1 INVX1_3013 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_3_), .Y(_20237_) );
	OAI21X1 OAI21X1_4473 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf87), .Y(_20238_) );
	AOI21X1 AOI21X1_2958 ( .gnd(gnd), .vdd(vdd), .A(_20237_), .B(_20231__bF_buf0), .C(_20238_), .Y(_17366__3_) );
	INVX1 INVX1_3014 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_4_), .Y(_20239_) );
	OAI21X1 OAI21X1_4474 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf86), .Y(_20240_) );
	AOI21X1 AOI21X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_20239_), .B(_20231__bF_buf6), .C(_20240_), .Y(_17366__4_) );
	INVX1 INVX1_3015 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_5_), .Y(_20241_) );
	OAI21X1 OAI21X1_4475 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf85), .Y(_20242_) );
	AOI21X1 AOI21X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_20241_), .B(_20231__bF_buf4), .C(_20242_), .Y(_17366__5_) );
	INVX1 INVX1_3016 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_6_), .Y(_20243_) );
	OAI21X1 OAI21X1_4476 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf84), .Y(_20244_) );
	AOI21X1 AOI21X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_20243_), .B(_20231__bF_buf2), .C(_20244_), .Y(_17366__6_) );
	INVX1 INVX1_3017 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_7_), .Y(_20245_) );
	OAI21X1 OAI21X1_4477 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf83), .Y(_20246_) );
	AOI21X1 AOI21X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_20245_), .B(_20231__bF_buf0), .C(_20246_), .Y(_17366__7_) );
	INVX1 INVX1_3018 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_8_), .Y(_20247_) );
	OAI21X1 OAI21X1_4478 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf82), .Y(_20248_) );
	AOI21X1 AOI21X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_20247_), .B(_20231__bF_buf6), .C(_20248_), .Y(_17366__8_) );
	INVX1 INVX1_3019 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_9_), .Y(_20249_) );
	OAI21X1 OAI21X1_4479 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf81), .Y(_20250_) );
	AOI21X1 AOI21X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_20249_), .B(_20231__bF_buf4), .C(_20250_), .Y(_17366__9_) );
	INVX1 INVX1_3020 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_10_), .Y(_20251_) );
	OAI21X1 OAI21X1_4480 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf80), .Y(_20252_) );
	AOI21X1 AOI21X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_20251_), .B(_20231__bF_buf2), .C(_20252_), .Y(_17366__10_) );
	INVX1 INVX1_3021 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_11_), .Y(_20253_) );
	OAI21X1 OAI21X1_4481 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf79), .Y(_20254_) );
	AOI21X1 AOI21X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_20253_), .B(_20231__bF_buf0), .C(_20254_), .Y(_17366__11_) );
	INVX1 INVX1_3022 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_12_), .Y(_20255_) );
	OAI21X1 OAI21X1_4482 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf78), .Y(_20256_) );
	AOI21X1 AOI21X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_20255_), .B(_20231__bF_buf6), .C(_20256_), .Y(_17366__12_) );
	INVX1 INVX1_3023 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_13_), .Y(_20257_) );
	OAI21X1 OAI21X1_4483 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf77), .Y(_20258_) );
	AOI21X1 AOI21X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_20257_), .B(_20231__bF_buf4), .C(_20258_), .Y(_17366__13_) );
	INVX1 INVX1_3024 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_14_), .Y(_20259_) );
	OAI21X1 OAI21X1_4484 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf76), .Y(_20260_) );
	AOI21X1 AOI21X1_2969 ( .gnd(gnd), .vdd(vdd), .A(_20259_), .B(_20231__bF_buf2), .C(_20260_), .Y(_17366__14_) );
	INVX1 INVX1_3025 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_15_), .Y(_20261_) );
	OAI21X1 OAI21X1_4485 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf75), .Y(_20262_) );
	AOI21X1 AOI21X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_20261_), .B(_20231__bF_buf0), .C(_20262_), .Y(_17366__15_) );
	INVX1 INVX1_3026 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_16_), .Y(_20263_) );
	OAI21X1 OAI21X1_4486 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf74), .Y(_20264_) );
	AOI21X1 AOI21X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_20263_), .B(_20231__bF_buf6), .C(_20264_), .Y(_17366__16_) );
	INVX1 INVX1_3027 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_17_), .Y(_20265_) );
	OAI21X1 OAI21X1_4487 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf73), .Y(_20266_) );
	AOI21X1 AOI21X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_20265_), .B(_20231__bF_buf4), .C(_20266_), .Y(_17366__17_) );
	INVX1 INVX1_3028 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_18_), .Y(_20267_) );
	OAI21X1 OAI21X1_4488 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf72), .Y(_20268_) );
	AOI21X1 AOI21X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_20267_), .B(_20231__bF_buf2), .C(_20268_), .Y(_17366__18_) );
	INVX1 INVX1_3029 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_19_), .Y(_20269_) );
	OAI21X1 OAI21X1_4489 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf71), .Y(_20270_) );
	AOI21X1 AOI21X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_20269_), .B(_20231__bF_buf0), .C(_20270_), .Y(_17366__19_) );
	INVX1 INVX1_3030 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_20_), .Y(_20271_) );
	OAI21X1 OAI21X1_4490 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf70), .Y(_20272_) );
	AOI21X1 AOI21X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_20271_), .B(_20231__bF_buf6), .C(_20272_), .Y(_17366__20_) );
	INVX1 INVX1_3031 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_21_), .Y(_20273_) );
	OAI21X1 OAI21X1_4491 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf69), .Y(_20274_) );
	AOI21X1 AOI21X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_20273_), .B(_20231__bF_buf4), .C(_20274_), .Y(_17366__21_) );
	INVX1 INVX1_3032 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_22_), .Y(_20275_) );
	OAI21X1 OAI21X1_4492 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf68), .Y(_20276_) );
	AOI21X1 AOI21X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_20275_), .B(_20231__bF_buf2), .C(_20276_), .Y(_17366__22_) );
	INVX1 INVX1_3033 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_23_), .Y(_20277_) );
	OAI21X1 OAI21X1_4493 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf67), .Y(_20278_) );
	AOI21X1 AOI21X1_2978 ( .gnd(gnd), .vdd(vdd), .A(_20277_), .B(_20231__bF_buf0), .C(_20278_), .Y(_17366__23_) );
	INVX1 INVX1_3034 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_24_), .Y(_20279_) );
	OAI21X1 OAI21X1_4494 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf66), .Y(_20280_) );
	AOI21X1 AOI21X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_20279_), .B(_20231__bF_buf6), .C(_20280_), .Y(_17366__24_) );
	INVX1 INVX1_3035 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_25_), .Y(_20281_) );
	OAI21X1 OAI21X1_4495 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf65), .Y(_20282_) );
	AOI21X1 AOI21X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_20281_), .B(_20231__bF_buf4), .C(_20282_), .Y(_17366__25_) );
	INVX1 INVX1_3036 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_26_), .Y(_20283_) );
	OAI21X1 OAI21X1_4496 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf64), .Y(_20284_) );
	AOI21X1 AOI21X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_20283_), .B(_20231__bF_buf2), .C(_20284_), .Y(_17366__26_) );
	INVX1 INVX1_3037 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_27_), .Y(_20285_) );
	OAI21X1 OAI21X1_4497 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf63), .Y(_20286_) );
	AOI21X1 AOI21X1_2982 ( .gnd(gnd), .vdd(vdd), .A(_20285_), .B(_20231__bF_buf0), .C(_20286_), .Y(_17366__27_) );
	INVX1 INVX1_3038 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_28_), .Y(_20287_) );
	OAI21X1 OAI21X1_4498 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_20231__bF_buf7), .C(_19153__bF_buf62), .Y(_20288_) );
	AOI21X1 AOI21X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_20287_), .B(_20231__bF_buf6), .C(_20288_), .Y(_17366__28_) );
	INVX1 INVX1_3039 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_29_), .Y(_20289_) );
	OAI21X1 OAI21X1_4499 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_20231__bF_buf5), .C(_19153__bF_buf61), .Y(_20290_) );
	AOI21X1 AOI21X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_20289_), .B(_20231__bF_buf4), .C(_20290_), .Y(_17366__29_) );
	INVX1 INVX1_3040 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_30_), .Y(_20291_) );
	OAI21X1 OAI21X1_4500 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_20231__bF_buf3), .C(_19153__bF_buf60), .Y(_20292_) );
	AOI21X1 AOI21X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_20291_), .B(_20231__bF_buf2), .C(_20292_), .Y(_17366__30_) );
	INVX1 INVX1_3041 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_31_), .Y(_20293_) );
	OAI21X1 OAI21X1_4501 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_20231__bF_buf1), .C(_19153__bF_buf59), .Y(_20294_) );
	AOI21X1 AOI21X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_20293_), .B(_20231__bF_buf0), .C(_20294_), .Y(_17366__31_) );
	INVX1 INVX1_3042 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_0_), .Y(_20295_) );
	NAND2X1 NAND2X1_3569 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19566_), .Y(_20296_) );
	OAI21X1 OAI21X1_4502 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf58), .Y(_20297_) );
	AOI21X1 AOI21X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_20295_), .B(_20296__bF_buf6), .C(_20297_), .Y(_17365__0_) );
	INVX1 INVX1_3043 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_1_), .Y(_20298_) );
	OAI21X1 OAI21X1_4503 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf57), .Y(_20299_) );
	AOI21X1 AOI21X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_20298_), .B(_20296__bF_buf4), .C(_20299_), .Y(_17365__1_) );
	INVX1 INVX1_3044 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_2_), .Y(_20300_) );
	OAI21X1 OAI21X1_4504 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf56), .Y(_20301_) );
	AOI21X1 AOI21X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_20300_), .B(_20296__bF_buf2), .C(_20301_), .Y(_17365__2_) );
	INVX1 INVX1_3045 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_3_), .Y(_20302_) );
	OAI21X1 OAI21X1_4505 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf55), .Y(_20303_) );
	AOI21X1 AOI21X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_20302_), .B(_20296__bF_buf0), .C(_20303_), .Y(_17365__3_) );
	INVX1 INVX1_3046 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_4_), .Y(_20304_) );
	OAI21X1 OAI21X1_4506 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf54), .Y(_20305_) );
	AOI21X1 AOI21X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_20304_), .B(_20296__bF_buf6), .C(_20305_), .Y(_17365__4_) );
	INVX1 INVX1_3047 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_5_), .Y(_20306_) );
	OAI21X1 OAI21X1_4507 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf53), .Y(_20307_) );
	AOI21X1 AOI21X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_20306_), .B(_20296__bF_buf4), .C(_20307_), .Y(_17365__5_) );
	INVX1 INVX1_3048 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_6_), .Y(_20308_) );
	OAI21X1 OAI21X1_4508 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf52), .Y(_20309_) );
	AOI21X1 AOI21X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_20308_), .B(_20296__bF_buf2), .C(_20309_), .Y(_17365__6_) );
	INVX1 INVX1_3049 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_7_), .Y(_20310_) );
	OAI21X1 OAI21X1_4509 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf51), .Y(_20311_) );
	AOI21X1 AOI21X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_20310_), .B(_20296__bF_buf0), .C(_20311_), .Y(_17365__7_) );
	INVX1 INVX1_3050 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_8_), .Y(_20312_) );
	OAI21X1 OAI21X1_4510 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf50), .Y(_20313_) );
	AOI21X1 AOI21X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_20312_), .B(_20296__bF_buf6), .C(_20313_), .Y(_17365__8_) );
	INVX1 INVX1_3051 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_9_), .Y(_20314_) );
	OAI21X1 OAI21X1_4511 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf49), .Y(_20315_) );
	AOI21X1 AOI21X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_20314_), .B(_20296__bF_buf4), .C(_20315_), .Y(_17365__9_) );
	INVX1 INVX1_3052 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_10_), .Y(_20316_) );
	OAI21X1 OAI21X1_4512 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf48), .Y(_20317_) );
	AOI21X1 AOI21X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_20316_), .B(_20296__bF_buf2), .C(_20317_), .Y(_17365__10_) );
	INVX1 INVX1_3053 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_11_), .Y(_20318_) );
	OAI21X1 OAI21X1_4513 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf47), .Y(_20319_) );
	AOI21X1 AOI21X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_20318_), .B(_20296__bF_buf0), .C(_20319_), .Y(_17365__11_) );
	INVX1 INVX1_3054 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_12_), .Y(_20320_) );
	OAI21X1 OAI21X1_4514 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf46), .Y(_20321_) );
	AOI21X1 AOI21X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_20320_), .B(_20296__bF_buf6), .C(_20321_), .Y(_17365__12_) );
	INVX1 INVX1_3055 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_13_), .Y(_20322_) );
	OAI21X1 OAI21X1_4515 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf45), .Y(_20323_) );
	AOI21X1 AOI21X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_20322_), .B(_20296__bF_buf4), .C(_20323_), .Y(_17365__13_) );
	INVX1 INVX1_3056 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_14_), .Y(_20324_) );
	OAI21X1 OAI21X1_4516 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf44), .Y(_20325_) );
	AOI21X1 AOI21X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_20324_), .B(_20296__bF_buf2), .C(_20325_), .Y(_17365__14_) );
	INVX1 INVX1_3057 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_15_), .Y(_20326_) );
	OAI21X1 OAI21X1_4517 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf43), .Y(_20327_) );
	AOI21X1 AOI21X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_20326_), .B(_20296__bF_buf0), .C(_20327_), .Y(_17365__15_) );
	INVX1 INVX1_3058 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_16_), .Y(_20328_) );
	OAI21X1 OAI21X1_4518 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf42), .Y(_20329_) );
	AOI21X1 AOI21X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_20328_), .B(_20296__bF_buf6), .C(_20329_), .Y(_17365__16_) );
	INVX1 INVX1_3059 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_17_), .Y(_20330_) );
	OAI21X1 OAI21X1_4519 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf41), .Y(_20331_) );
	AOI21X1 AOI21X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_20330_), .B(_20296__bF_buf4), .C(_20331_), .Y(_17365__17_) );
	INVX1 INVX1_3060 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_18_), .Y(_20332_) );
	OAI21X1 OAI21X1_4520 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf40), .Y(_20333_) );
	AOI21X1 AOI21X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_20332_), .B(_20296__bF_buf2), .C(_20333_), .Y(_17365__18_) );
	INVX1 INVX1_3061 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_19_), .Y(_20334_) );
	OAI21X1 OAI21X1_4521 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf39), .Y(_20335_) );
	AOI21X1 AOI21X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_20334_), .B(_20296__bF_buf0), .C(_20335_), .Y(_17365__19_) );
	INVX1 INVX1_3062 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_20_), .Y(_20336_) );
	OAI21X1 OAI21X1_4522 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf38), .Y(_20337_) );
	AOI21X1 AOI21X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_20336_), .B(_20296__bF_buf6), .C(_20337_), .Y(_17365__20_) );
	INVX1 INVX1_3063 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_21_), .Y(_20338_) );
	OAI21X1 OAI21X1_4523 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf37), .Y(_20339_) );
	AOI21X1 AOI21X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_20338_), .B(_20296__bF_buf4), .C(_20339_), .Y(_17365__21_) );
	INVX1 INVX1_3064 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_22_), .Y(_20340_) );
	OAI21X1 OAI21X1_4524 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf36), .Y(_20341_) );
	AOI21X1 AOI21X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_20340_), .B(_20296__bF_buf2), .C(_20341_), .Y(_17365__22_) );
	INVX1 INVX1_3065 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_23_), .Y(_20342_) );
	OAI21X1 OAI21X1_4525 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf35), .Y(_20343_) );
	AOI21X1 AOI21X1_3010 ( .gnd(gnd), .vdd(vdd), .A(_20342_), .B(_20296__bF_buf0), .C(_20343_), .Y(_17365__23_) );
	INVX1 INVX1_3066 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_24_), .Y(_20344_) );
	OAI21X1 OAI21X1_4526 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf34), .Y(_20345_) );
	AOI21X1 AOI21X1_3011 ( .gnd(gnd), .vdd(vdd), .A(_20344_), .B(_20296__bF_buf6), .C(_20345_), .Y(_17365__24_) );
	INVX1 INVX1_3067 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_25_), .Y(_20346_) );
	OAI21X1 OAI21X1_4527 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf33), .Y(_20347_) );
	AOI21X1 AOI21X1_3012 ( .gnd(gnd), .vdd(vdd), .A(_20346_), .B(_20296__bF_buf4), .C(_20347_), .Y(_17365__25_) );
	INVX1 INVX1_3068 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_26_), .Y(_20348_) );
	OAI21X1 OAI21X1_4528 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf32), .Y(_20349_) );
	AOI21X1 AOI21X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_20348_), .B(_20296__bF_buf2), .C(_20349_), .Y(_17365__26_) );
	INVX1 INVX1_3069 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_27_), .Y(_20350_) );
	OAI21X1 OAI21X1_4529 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf31), .Y(_20351_) );
	AOI21X1 AOI21X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_20350_), .B(_20296__bF_buf0), .C(_20351_), .Y(_17365__27_) );
	INVX1 INVX1_3070 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_28_), .Y(_20352_) );
	OAI21X1 OAI21X1_4530 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf3), .B(_20296__bF_buf7), .C(_19153__bF_buf30), .Y(_20353_) );
	AOI21X1 AOI21X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_20352_), .B(_20296__bF_buf6), .C(_20353_), .Y(_17365__28_) );
	INVX1 INVX1_3071 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_29_), .Y(_20354_) );
	OAI21X1 OAI21X1_4531 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf3), .B(_20296__bF_buf5), .C(_19153__bF_buf29), .Y(_20355_) );
	AOI21X1 AOI21X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_20354_), .B(_20296__bF_buf4), .C(_20355_), .Y(_17365__29_) );
	INVX1 INVX1_3072 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_30_), .Y(_20356_) );
	OAI21X1 OAI21X1_4532 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf3), .B(_20296__bF_buf3), .C(_19153__bF_buf28), .Y(_20357_) );
	AOI21X1 AOI21X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_20356_), .B(_20296__bF_buf2), .C(_20357_), .Y(_17365__30_) );
	INVX1 INVX1_3073 ( .gnd(gnd), .vdd(vdd), .A(registers_r5_31_), .Y(_20358_) );
	OAI21X1 OAI21X1_4533 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf3), .B(_20296__bF_buf1), .C(_19153__bF_buf27), .Y(_20359_) );
	AOI21X1 AOI21X1_3018 ( .gnd(gnd), .vdd(vdd), .A(_20358_), .B(_20296__bF_buf0), .C(_20359_), .Y(_17365__31_) );
	INVX1 INVX1_3074 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_0_), .Y(_20360_) );
	NAND2X1 NAND2X1_3570 ( .gnd(gnd), .vdd(vdd), .A(_19601_), .B(_20100_), .Y(_20361_) );
	OAI21X1 OAI21X1_4534 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf26), .Y(_20362_) );
	AOI21X1 AOI21X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_20360_), .B(_20361__bF_buf6), .C(_20362_), .Y(_17364__0_) );
	INVX1 INVX1_3075 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_1_), .Y(_20363_) );
	OAI21X1 OAI21X1_4535 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf25), .Y(_20364_) );
	AOI21X1 AOI21X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_20363_), .B(_20361__bF_buf4), .C(_20364_), .Y(_17364__1_) );
	INVX1 INVX1_3076 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_2_), .Y(_20365_) );
	OAI21X1 OAI21X1_4536 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf24), .Y(_20366_) );
	AOI21X1 AOI21X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_20365_), .B(_20361__bF_buf2), .C(_20366_), .Y(_17364__2_) );
	INVX1 INVX1_3077 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_3_), .Y(_20367_) );
	OAI21X1 OAI21X1_4537 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf23), .Y(_20368_) );
	AOI21X1 AOI21X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_20367_), .B(_20361__bF_buf0), .C(_20368_), .Y(_17364__3_) );
	INVX1 INVX1_3078 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_4_), .Y(_20369_) );
	OAI21X1 OAI21X1_4538 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf22), .Y(_20370_) );
	AOI21X1 AOI21X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_20369_), .B(_20361__bF_buf6), .C(_20370_), .Y(_17364__4_) );
	INVX1 INVX1_3079 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_5_), .Y(_20371_) );
	OAI21X1 OAI21X1_4539 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf21), .Y(_20372_) );
	AOI21X1 AOI21X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_20371_), .B(_20361__bF_buf4), .C(_20372_), .Y(_17364__5_) );
	INVX1 INVX1_3080 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_6_), .Y(_20373_) );
	OAI21X1 OAI21X1_4540 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf20), .Y(_20374_) );
	AOI21X1 AOI21X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_20373_), .B(_20361__bF_buf2), .C(_20374_), .Y(_17364__6_) );
	INVX1 INVX1_3081 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_7_), .Y(_20375_) );
	OAI21X1 OAI21X1_4541 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf19), .Y(_20376_) );
	AOI21X1 AOI21X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_20375_), .B(_20361__bF_buf0), .C(_20376_), .Y(_17364__7_) );
	INVX1 INVX1_3082 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_8_), .Y(_20377_) );
	OAI21X1 OAI21X1_4542 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf18), .Y(_20378_) );
	AOI21X1 AOI21X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_20377_), .B(_20361__bF_buf6), .C(_20378_), .Y(_17364__8_) );
	INVX1 INVX1_3083 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_9_), .Y(_20379_) );
	OAI21X1 OAI21X1_4543 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf17), .Y(_20380_) );
	AOI21X1 AOI21X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_20379_), .B(_20361__bF_buf4), .C(_20380_), .Y(_17364__9_) );
	INVX1 INVX1_3084 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_10_), .Y(_20381_) );
	OAI21X1 OAI21X1_4544 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf16), .Y(_20382_) );
	AOI21X1 AOI21X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_20381_), .B(_20361__bF_buf2), .C(_20382_), .Y(_17364__10_) );
	INVX1 INVX1_3085 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_11_), .Y(_20383_) );
	OAI21X1 OAI21X1_4545 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf15), .Y(_20384_) );
	AOI21X1 AOI21X1_3030 ( .gnd(gnd), .vdd(vdd), .A(_20383_), .B(_20361__bF_buf0), .C(_20384_), .Y(_17364__11_) );
	INVX1 INVX1_3086 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_12_), .Y(_20385_) );
	OAI21X1 OAI21X1_4546 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf14), .Y(_20386_) );
	AOI21X1 AOI21X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_20385_), .B(_20361__bF_buf6), .C(_20386_), .Y(_17364__12_) );
	INVX1 INVX1_3087 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_13_), .Y(_20387_) );
	OAI21X1 OAI21X1_4547 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf13), .Y(_20388_) );
	AOI21X1 AOI21X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_20387_), .B(_20361__bF_buf4), .C(_20388_), .Y(_17364__13_) );
	INVX1 INVX1_3088 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_14_), .Y(_20389_) );
	OAI21X1 OAI21X1_4548 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf12), .Y(_20390_) );
	AOI21X1 AOI21X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_20389_), .B(_20361__bF_buf2), .C(_20390_), .Y(_17364__14_) );
	INVX1 INVX1_3089 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_15_), .Y(_20391_) );
	OAI21X1 OAI21X1_4549 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf11), .Y(_20392_) );
	AOI21X1 AOI21X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_20391_), .B(_20361__bF_buf0), .C(_20392_), .Y(_17364__15_) );
	INVX1 INVX1_3090 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_16_), .Y(_20393_) );
	OAI21X1 OAI21X1_4550 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf10), .Y(_20394_) );
	AOI21X1 AOI21X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_20393_), .B(_20361__bF_buf6), .C(_20394_), .Y(_17364__16_) );
	INVX1 INVX1_3091 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_17_), .Y(_20395_) );
	OAI21X1 OAI21X1_4551 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf9), .Y(_20396_) );
	AOI21X1 AOI21X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_20395_), .B(_20361__bF_buf4), .C(_20396_), .Y(_17364__17_) );
	INVX1 INVX1_3092 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_18_), .Y(_20397_) );
	OAI21X1 OAI21X1_4552 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf8), .Y(_20398_) );
	AOI21X1 AOI21X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_20397_), .B(_20361__bF_buf2), .C(_20398_), .Y(_17364__18_) );
	INVX1 INVX1_3093 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_19_), .Y(_20399_) );
	OAI21X1 OAI21X1_4553 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf7), .Y(_20400_) );
	AOI21X1 AOI21X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_20399_), .B(_20361__bF_buf0), .C(_20400_), .Y(_17364__19_) );
	INVX1 INVX1_3094 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_20_), .Y(_20401_) );
	OAI21X1 OAI21X1_4554 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf6), .Y(_20402_) );
	AOI21X1 AOI21X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_20401_), .B(_20361__bF_buf6), .C(_20402_), .Y(_17364__20_) );
	INVX1 INVX1_3095 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_21_), .Y(_20403_) );
	OAI21X1 OAI21X1_4555 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf5), .Y(_20404_) );
	AOI21X1 AOI21X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_20403_), .B(_20361__bF_buf4), .C(_20404_), .Y(_17364__21_) );
	INVX1 INVX1_3096 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_22_), .Y(_20405_) );
	OAI21X1 OAI21X1_4556 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf4), .Y(_20406_) );
	AOI21X1 AOI21X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_20405_), .B(_20361__bF_buf2), .C(_20406_), .Y(_17364__22_) );
	INVX1 INVX1_3097 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_23_), .Y(_20407_) );
	OAI21X1 OAI21X1_4557 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf3), .Y(_20408_) );
	AOI21X1 AOI21X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_20407_), .B(_20361__bF_buf0), .C(_20408_), .Y(_17364__23_) );
	INVX1 INVX1_3098 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_24_), .Y(_20409_) );
	OAI21X1 OAI21X1_4558 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf2), .Y(_20410_) );
	AOI21X1 AOI21X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_20409_), .B(_20361__bF_buf6), .C(_20410_), .Y(_17364__24_) );
	INVX1 INVX1_3099 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_25_), .Y(_20411_) );
	OAI21X1 OAI21X1_4559 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf1), .Y(_20412_) );
	AOI21X1 AOI21X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_20411_), .B(_20361__bF_buf4), .C(_20412_), .Y(_17364__25_) );
	INVX1 INVX1_3100 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_26_), .Y(_20413_) );
	OAI21X1 OAI21X1_4560 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf0), .Y(_20414_) );
	AOI21X1 AOI21X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_20413_), .B(_20361__bF_buf2), .C(_20414_), .Y(_17364__26_) );
	INVX1 INVX1_3101 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_27_), .Y(_20415_) );
	OAI21X1 OAI21X1_4561 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf98), .Y(_20416_) );
	AOI21X1 AOI21X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_20415_), .B(_20361__bF_buf0), .C(_20416_), .Y(_17364__27_) );
	INVX1 INVX1_3102 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_28_), .Y(_20417_) );
	OAI21X1 OAI21X1_4562 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf2), .B(_20361__bF_buf7), .C(_19153__bF_buf97), .Y(_20418_) );
	AOI21X1 AOI21X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_20417_), .B(_20361__bF_buf6), .C(_20418_), .Y(_17364__28_) );
	INVX1 INVX1_3103 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_29_), .Y(_20419_) );
	OAI21X1 OAI21X1_4563 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf2), .B(_20361__bF_buf5), .C(_19153__bF_buf96), .Y(_20420_) );
	AOI21X1 AOI21X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_20419_), .B(_20361__bF_buf4), .C(_20420_), .Y(_17364__29_) );
	INVX1 INVX1_3104 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_30_), .Y(_20421_) );
	OAI21X1 OAI21X1_4564 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf2), .B(_20361__bF_buf3), .C(_19153__bF_buf95), .Y(_20422_) );
	AOI21X1 AOI21X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_20421_), .B(_20361__bF_buf2), .C(_20422_), .Y(_17364__30_) );
	INVX1 INVX1_3105 ( .gnd(gnd), .vdd(vdd), .A(registers_r4_31_), .Y(_20423_) );
	OAI21X1 OAI21X1_4565 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf2), .B(_20361__bF_buf1), .C(_19153__bF_buf94), .Y(_20424_) );
	AOI21X1 AOI21X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_20423_), .B(_20361__bF_buf0), .C(_20424_), .Y(_17364__31_) );
	NAND2X1 NAND2X1_3571 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19667_), .Y(_20425_) );
	OAI21X1 OAI21X1_4566 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf93), .Y(_20426_) );
	AOI21X1 AOI21X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_17379_), .B(_20425__bF_buf6), .C(_20426_), .Y(_17363__0_) );
	OAI21X1 OAI21X1_4567 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf92), .Y(_20427_) );
	AOI21X1 AOI21X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_17475_), .B(_20425__bF_buf4), .C(_20427_), .Y(_17363__1_) );
	OAI21X1 OAI21X1_4568 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf91), .Y(_20428_) );
	AOI21X1 AOI21X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_17529_), .B(_20425__bF_buf2), .C(_20428_), .Y(_17363__2_) );
	OAI21X1 OAI21X1_4569 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf90), .Y(_20429_) );
	AOI21X1 AOI21X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_17583_), .B(_20425__bF_buf0), .C(_20429_), .Y(_17363__3_) );
	OAI21X1 OAI21X1_4570 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf89), .Y(_20430_) );
	AOI21X1 AOI21X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_17637_), .B(_20425__bF_buf6), .C(_20430_), .Y(_17363__4_) );
	OAI21X1 OAI21X1_4571 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf88), .Y(_20431_) );
	AOI21X1 AOI21X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_17691_), .B(_20425__bF_buf4), .C(_20431_), .Y(_17363__5_) );
	OAI21X1 OAI21X1_4572 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf87), .Y(_20432_) );
	AOI21X1 AOI21X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_17745_), .B(_20425__bF_buf2), .C(_20432_), .Y(_17363__6_) );
	OAI21X1 OAI21X1_4573 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf86), .Y(_20433_) );
	AOI21X1 AOI21X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_17799_), .B(_20425__bF_buf0), .C(_20433_), .Y(_17363__7_) );
	OAI21X1 OAI21X1_4574 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf85), .Y(_20434_) );
	AOI21X1 AOI21X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_17853_), .B(_20425__bF_buf6), .C(_20434_), .Y(_17363__8_) );
	OAI21X1 OAI21X1_4575 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf84), .Y(_20435_) );
	AOI21X1 AOI21X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_17907_), .B(_20425__bF_buf4), .C(_20435_), .Y(_17363__9_) );
	OAI21X1 OAI21X1_4576 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf83), .Y(_20436_) );
	AOI21X1 AOI21X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_17961_), .B(_20425__bF_buf2), .C(_20436_), .Y(_17363__10_) );
	OAI21X1 OAI21X1_4577 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf82), .Y(_20437_) );
	AOI21X1 AOI21X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_18015_), .B(_20425__bF_buf0), .C(_20437_), .Y(_17363__11_) );
	OAI21X1 OAI21X1_4578 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf81), .Y(_20438_) );
	AOI21X1 AOI21X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_18069_), .B(_20425__bF_buf6), .C(_20438_), .Y(_17363__12_) );
	OAI21X1 OAI21X1_4579 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf80), .Y(_20439_) );
	AOI21X1 AOI21X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_18123_), .B(_20425__bF_buf4), .C(_20439_), .Y(_17363__13_) );
	OAI21X1 OAI21X1_4580 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf79), .Y(_20440_) );
	AOI21X1 AOI21X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_18177_), .B(_20425__bF_buf2), .C(_20440_), .Y(_17363__14_) );
	OAI21X1 OAI21X1_4581 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf78), .Y(_20441_) );
	AOI21X1 AOI21X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_18231_), .B(_20425__bF_buf0), .C(_20441_), .Y(_17363__15_) );
	OAI21X1 OAI21X1_4582 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf77), .Y(_20442_) );
	AOI21X1 AOI21X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_18285_), .B(_20425__bF_buf6), .C(_20442_), .Y(_17363__16_) );
	OAI21X1 OAI21X1_4583 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf76), .Y(_20443_) );
	AOI21X1 AOI21X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_18339_), .B(_20425__bF_buf4), .C(_20443_), .Y(_17363__17_) );
	OAI21X1 OAI21X1_4584 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf75), .Y(_20444_) );
	AOI21X1 AOI21X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_18393_), .B(_20425__bF_buf2), .C(_20444_), .Y(_17363__18_) );
	OAI21X1 OAI21X1_4585 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf74), .Y(_20445_) );
	AOI21X1 AOI21X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_18447_), .B(_20425__bF_buf0), .C(_20445_), .Y(_17363__19_) );
	OAI21X1 OAI21X1_4586 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf73), .Y(_20446_) );
	AOI21X1 AOI21X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_18501_), .B(_20425__bF_buf6), .C(_20446_), .Y(_17363__20_) );
	OAI21X1 OAI21X1_4587 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf72), .Y(_20447_) );
	AOI21X1 AOI21X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_18555_), .B(_20425__bF_buf4), .C(_20447_), .Y(_17363__21_) );
	OAI21X1 OAI21X1_4588 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf71), .Y(_20448_) );
	AOI21X1 AOI21X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_18609_), .B(_20425__bF_buf2), .C(_20448_), .Y(_17363__22_) );
	OAI21X1 OAI21X1_4589 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf70), .Y(_20449_) );
	AOI21X1 AOI21X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_18663_), .B(_20425__bF_buf0), .C(_20449_), .Y(_17363__23_) );
	OAI21X1 OAI21X1_4590 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf69), .Y(_20450_) );
	AOI21X1 AOI21X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_18717_), .B(_20425__bF_buf6), .C(_20450_), .Y(_17363__24_) );
	OAI21X1 OAI21X1_4591 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf68), .Y(_20451_) );
	AOI21X1 AOI21X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_18771_), .B(_20425__bF_buf4), .C(_20451_), .Y(_17363__25_) );
	OAI21X1 OAI21X1_4592 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf67), .Y(_20452_) );
	AOI21X1 AOI21X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_18825_), .B(_20425__bF_buf2), .C(_20452_), .Y(_17363__26_) );
	OAI21X1 OAI21X1_4593 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf66), .Y(_20453_) );
	AOI21X1 AOI21X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_18879_), .B(_20425__bF_buf0), .C(_20453_), .Y(_17363__27_) );
	OAI21X1 OAI21X1_4594 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf1), .B(_20425__bF_buf7), .C(_19153__bF_buf65), .Y(_20454_) );
	AOI21X1 AOI21X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_18933_), .B(_20425__bF_buf6), .C(_20454_), .Y(_17363__28_) );
	OAI21X1 OAI21X1_4595 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf1), .B(_20425__bF_buf5), .C(_19153__bF_buf64), .Y(_20455_) );
	AOI21X1 AOI21X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_18987_), .B(_20425__bF_buf4), .C(_20455_), .Y(_17363__29_) );
	OAI21X1 OAI21X1_4596 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf1), .B(_20425__bF_buf3), .C(_19153__bF_buf63), .Y(_20456_) );
	AOI21X1 AOI21X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_19041_), .B(_20425__bF_buf2), .C(_20456_), .Y(_17363__30_) );
	OAI21X1 OAI21X1_4597 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf1), .B(_20425__bF_buf1), .C(_19153__bF_buf62), .Y(_20457_) );
	AOI21X1 AOI21X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_19095_), .B(_20425__bF_buf0), .C(_20457_), .Y(_17363__31_) );
	NAND2X1 NAND2X1_3572 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19701_), .Y(_20458_) );
	OAI21X1 OAI21X1_4598 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf61), .Y(_20459_) );
	AOI21X1 AOI21X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_17380_), .B(_20458__bF_buf6), .C(_20459_), .Y(_17360__0_) );
	OAI21X1 OAI21X1_4599 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf60), .Y(_20460_) );
	AOI21X1 AOI21X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_17476_), .B(_20458__bF_buf4), .C(_20460_), .Y(_17360__1_) );
	OAI21X1 OAI21X1_4600 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf59), .Y(_20461_) );
	AOI21X1 AOI21X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_17530_), .B(_20458__bF_buf2), .C(_20461_), .Y(_17360__2_) );
	OAI21X1 OAI21X1_4601 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf58), .Y(_20462_) );
	AOI21X1 AOI21X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_17584_), .B(_20458__bF_buf0), .C(_20462_), .Y(_17360__3_) );
	OAI21X1 OAI21X1_4602 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf57), .Y(_20463_) );
	AOI21X1 AOI21X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_17638_), .B(_20458__bF_buf6), .C(_20463_), .Y(_17360__4_) );
	OAI21X1 OAI21X1_4603 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf56), .Y(_20464_) );
	AOI21X1 AOI21X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_17692_), .B(_20458__bF_buf4), .C(_20464_), .Y(_17360__5_) );
	OAI21X1 OAI21X1_4604 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf55), .Y(_20465_) );
	AOI21X1 AOI21X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_17746_), .B(_20458__bF_buf2), .C(_20465_), .Y(_17360__6_) );
	OAI21X1 OAI21X1_4605 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf54), .Y(_20466_) );
	AOI21X1 AOI21X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_17800_), .B(_20458__bF_buf0), .C(_20466_), .Y(_17360__7_) );
	OAI21X1 OAI21X1_4606 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf53), .Y(_20467_) );
	AOI21X1 AOI21X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_17854_), .B(_20458__bF_buf6), .C(_20467_), .Y(_17360__8_) );
	OAI21X1 OAI21X1_4607 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf52), .Y(_20468_) );
	AOI21X1 AOI21X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_17908_), .B(_20458__bF_buf4), .C(_20468_), .Y(_17360__9_) );
	OAI21X1 OAI21X1_4608 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf51), .Y(_20469_) );
	AOI21X1 AOI21X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_17962_), .B(_20458__bF_buf2), .C(_20469_), .Y(_17360__10_) );
	OAI21X1 OAI21X1_4609 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf50), .Y(_20470_) );
	AOI21X1 AOI21X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_18016_), .B(_20458__bF_buf0), .C(_20470_), .Y(_17360__11_) );
	OAI21X1 OAI21X1_4610 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf49), .Y(_20471_) );
	AOI21X1 AOI21X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_18070_), .B(_20458__bF_buf6), .C(_20471_), .Y(_17360__12_) );
	OAI21X1 OAI21X1_4611 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf48), .Y(_20472_) );
	AOI21X1 AOI21X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_18124_), .B(_20458__bF_buf4), .C(_20472_), .Y(_17360__13_) );
	OAI21X1 OAI21X1_4612 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf47), .Y(_20473_) );
	AOI21X1 AOI21X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_18178_), .B(_20458__bF_buf2), .C(_20473_), .Y(_17360__14_) );
	OAI21X1 OAI21X1_4613 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf46), .Y(_20474_) );
	AOI21X1 AOI21X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_18232_), .B(_20458__bF_buf0), .C(_20474_), .Y(_17360__15_) );
	OAI21X1 OAI21X1_4614 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf45), .Y(_20475_) );
	AOI21X1 AOI21X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_18286_), .B(_20458__bF_buf6), .C(_20475_), .Y(_17360__16_) );
	OAI21X1 OAI21X1_4615 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf44), .Y(_20476_) );
	AOI21X1 AOI21X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_18340_), .B(_20458__bF_buf4), .C(_20476_), .Y(_17360__17_) );
	OAI21X1 OAI21X1_4616 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf43), .Y(_20477_) );
	AOI21X1 AOI21X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_18394_), .B(_20458__bF_buf2), .C(_20477_), .Y(_17360__18_) );
	OAI21X1 OAI21X1_4617 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf42), .Y(_20478_) );
	AOI21X1 AOI21X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_18448_), .B(_20458__bF_buf0), .C(_20478_), .Y(_17360__19_) );
	OAI21X1 OAI21X1_4618 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf41), .Y(_20479_) );
	AOI21X1 AOI21X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_18502_), .B(_20458__bF_buf6), .C(_20479_), .Y(_17360__20_) );
	OAI21X1 OAI21X1_4619 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf40), .Y(_20480_) );
	AOI21X1 AOI21X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_18556_), .B(_20458__bF_buf4), .C(_20480_), .Y(_17360__21_) );
	OAI21X1 OAI21X1_4620 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf39), .Y(_20481_) );
	AOI21X1 AOI21X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_18610_), .B(_20458__bF_buf2), .C(_20481_), .Y(_17360__22_) );
	OAI21X1 OAI21X1_4621 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf38), .Y(_20482_) );
	AOI21X1 AOI21X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_18664_), .B(_20458__bF_buf0), .C(_20482_), .Y(_17360__23_) );
	OAI21X1 OAI21X1_4622 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf37), .Y(_20483_) );
	AOI21X1 AOI21X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_18718_), .B(_20458__bF_buf6), .C(_20483_), .Y(_17360__24_) );
	OAI21X1 OAI21X1_4623 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf36), .Y(_20484_) );
	AOI21X1 AOI21X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_18772_), .B(_20458__bF_buf4), .C(_20484_), .Y(_17360__25_) );
	OAI21X1 OAI21X1_4624 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf35), .Y(_20485_) );
	AOI21X1 AOI21X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_18826_), .B(_20458__bF_buf2), .C(_20485_), .Y(_17360__26_) );
	OAI21X1 OAI21X1_4625 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf34), .Y(_20486_) );
	AOI21X1 AOI21X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_18880_), .B(_20458__bF_buf0), .C(_20486_), .Y(_17360__27_) );
	OAI21X1 OAI21X1_4626 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf0), .B(_20458__bF_buf7), .C(_19153__bF_buf33), .Y(_20487_) );
	AOI21X1 AOI21X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_18934_), .B(_20458__bF_buf6), .C(_20487_), .Y(_17360__28_) );
	OAI21X1 OAI21X1_4627 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf0), .B(_20458__bF_buf5), .C(_19153__bF_buf32), .Y(_20488_) );
	AOI21X1 AOI21X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_18988_), .B(_20458__bF_buf4), .C(_20488_), .Y(_17360__29_) );
	OAI21X1 OAI21X1_4628 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf0), .B(_20458__bF_buf3), .C(_19153__bF_buf31), .Y(_20489_) );
	AOI21X1 AOI21X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_19042_), .B(_20458__bF_buf2), .C(_20489_), .Y(_17360__30_) );
	OAI21X1 OAI21X1_4629 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf0), .B(_20458__bF_buf1), .C(_19153__bF_buf30), .Y(_20490_) );
	AOI21X1 AOI21X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_19096_), .B(_20458__bF_buf0), .C(_20490_), .Y(_17360__31_) );
	INVX1 INVX1_3106 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_0_), .Y(_20491_) );
	NAND2X1 NAND2X1_3573 ( .gnd(gnd), .vdd(vdd), .A(_19803_), .B(_19735_), .Y(_20492_) );
	OAI21X1 OAI21X1_4630 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_0_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf29), .Y(_20493_) );
	AOI21X1 AOI21X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_20491_), .B(_20492__bF_buf6), .C(_20493_), .Y(_17349__0_) );
	INVX1 INVX1_3107 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_1_), .Y(_20494_) );
	OAI21X1 OAI21X1_4631 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_1_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf28), .Y(_20495_) );
	AOI21X1 AOI21X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_20494_), .B(_20492__bF_buf4), .C(_20495_), .Y(_17349__1_) );
	INVX1 INVX1_3108 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_2_), .Y(_20496_) );
	OAI21X1 OAI21X1_4632 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_2_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf27), .Y(_20497_) );
	AOI21X1 AOI21X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_20496_), .B(_20492__bF_buf2), .C(_20497_), .Y(_17349__2_) );
	INVX1 INVX1_3109 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_3_), .Y(_20498_) );
	OAI21X1 OAI21X1_4633 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_3_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf26), .Y(_20499_) );
	AOI21X1 AOI21X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_20498_), .B(_20492__bF_buf0), .C(_20499_), .Y(_17349__3_) );
	INVX1 INVX1_3110 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_4_), .Y(_20500_) );
	OAI21X1 OAI21X1_4634 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_4_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf25), .Y(_20501_) );
	AOI21X1 AOI21X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_20500_), .B(_20492__bF_buf6), .C(_20501_), .Y(_17349__4_) );
	INVX1 INVX1_3111 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_5_), .Y(_20502_) );
	OAI21X1 OAI21X1_4635 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_5_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf24), .Y(_20503_) );
	AOI21X1 AOI21X1_3120 ( .gnd(gnd), .vdd(vdd), .A(_20502_), .B(_20492__bF_buf4), .C(_20503_), .Y(_17349__5_) );
	INVX1 INVX1_3112 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_6_), .Y(_20504_) );
	OAI21X1 OAI21X1_4636 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_6_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf23), .Y(_20505_) );
	AOI21X1 AOI21X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_20504_), .B(_20492__bF_buf2), .C(_20505_), .Y(_17349__6_) );
	INVX1 INVX1_3113 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_7_), .Y(_20506_) );
	OAI21X1 OAI21X1_4637 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_7_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf22), .Y(_20507_) );
	AOI21X1 AOI21X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_20506_), .B(_20492__bF_buf0), .C(_20507_), .Y(_17349__7_) );
	INVX1 INVX1_3114 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_8_), .Y(_20508_) );
	OAI21X1 OAI21X1_4638 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_8_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf21), .Y(_20509_) );
	AOI21X1 AOI21X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_20508_), .B(_20492__bF_buf6), .C(_20509_), .Y(_17349__8_) );
	INVX1 INVX1_3115 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_9_), .Y(_20510_) );
	OAI21X1 OAI21X1_4639 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_9_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf20), .Y(_20511_) );
	AOI21X1 AOI21X1_3124 ( .gnd(gnd), .vdd(vdd), .A(_20510_), .B(_20492__bF_buf4), .C(_20511_), .Y(_17349__9_) );
	INVX1 INVX1_3116 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_10_), .Y(_20512_) );
	OAI21X1 OAI21X1_4640 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_10_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf19), .Y(_20513_) );
	AOI21X1 AOI21X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_20512_), .B(_20492__bF_buf2), .C(_20513_), .Y(_17349__10_) );
	INVX1 INVX1_3117 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_11_), .Y(_20514_) );
	OAI21X1 OAI21X1_4641 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_11_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf18), .Y(_20515_) );
	AOI21X1 AOI21X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_20514_), .B(_20492__bF_buf0), .C(_20515_), .Y(_17349__11_) );
	INVX1 INVX1_3118 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_12_), .Y(_20516_) );
	OAI21X1 OAI21X1_4642 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_12_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf17), .Y(_20517_) );
	AOI21X1 AOI21X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_20516_), .B(_20492__bF_buf6), .C(_20517_), .Y(_17349__12_) );
	INVX1 INVX1_3119 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_13_), .Y(_20518_) );
	OAI21X1 OAI21X1_4643 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_13_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf16), .Y(_20519_) );
	AOI21X1 AOI21X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_20518_), .B(_20492__bF_buf4), .C(_20519_), .Y(_17349__13_) );
	INVX1 INVX1_3120 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_14_), .Y(_20520_) );
	OAI21X1 OAI21X1_4644 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_14_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf15), .Y(_20521_) );
	AOI21X1 AOI21X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_20520_), .B(_20492__bF_buf2), .C(_20521_), .Y(_17349__14_) );
	INVX1 INVX1_3121 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_15_), .Y(_20522_) );
	OAI21X1 OAI21X1_4645 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_15_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf14), .Y(_20523_) );
	AOI21X1 AOI21X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_20522_), .B(_20492__bF_buf0), .C(_20523_), .Y(_17349__15_) );
	INVX1 INVX1_3122 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_16_), .Y(_20524_) );
	OAI21X1 OAI21X1_4646 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_16_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf13), .Y(_20525_) );
	AOI21X1 AOI21X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_20524_), .B(_20492__bF_buf6), .C(_20525_), .Y(_17349__16_) );
	INVX1 INVX1_3123 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_17_), .Y(_20526_) );
	OAI21X1 OAI21X1_4647 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_17_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf12), .Y(_20527_) );
	AOI21X1 AOI21X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_20526_), .B(_20492__bF_buf4), .C(_20527_), .Y(_17349__17_) );
	INVX1 INVX1_3124 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_18_), .Y(_20528_) );
	OAI21X1 OAI21X1_4648 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_18_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf11), .Y(_20529_) );
	AOI21X1 AOI21X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_20528_), .B(_20492__bF_buf2), .C(_20529_), .Y(_17349__18_) );
	INVX1 INVX1_3125 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_19_), .Y(_20530_) );
	OAI21X1 OAI21X1_4649 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_19_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf10), .Y(_20531_) );
	AOI21X1 AOI21X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_20530_), .B(_20492__bF_buf0), .C(_20531_), .Y(_17349__19_) );
	INVX1 INVX1_3126 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_20_), .Y(_20532_) );
	OAI21X1 OAI21X1_4650 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_20_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf9), .Y(_20533_) );
	AOI21X1 AOI21X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_20532_), .B(_20492__bF_buf6), .C(_20533_), .Y(_17349__20_) );
	INVX1 INVX1_3127 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_21_), .Y(_20534_) );
	OAI21X1 OAI21X1_4651 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_21_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf8), .Y(_20535_) );
	AOI21X1 AOI21X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_20534_), .B(_20492__bF_buf4), .C(_20535_), .Y(_17349__21_) );
	INVX1 INVX1_3128 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_22_), .Y(_20536_) );
	OAI21X1 OAI21X1_4652 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_22_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf7), .Y(_20537_) );
	AOI21X1 AOI21X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_20536_), .B(_20492__bF_buf2), .C(_20537_), .Y(_17349__22_) );
	INVX1 INVX1_3129 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_23_), .Y(_20538_) );
	OAI21X1 OAI21X1_4653 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_23_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf6), .Y(_20539_) );
	AOI21X1 AOI21X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_20538_), .B(_20492__bF_buf0), .C(_20539_), .Y(_17349__23_) );
	INVX1 INVX1_3130 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_24_), .Y(_20540_) );
	OAI21X1 OAI21X1_4654 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_24_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf5), .Y(_20541_) );
	AOI21X1 AOI21X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_20540_), .B(_20492__bF_buf6), .C(_20541_), .Y(_17349__24_) );
	INVX1 INVX1_3131 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_25_), .Y(_20542_) );
	OAI21X1 OAI21X1_4655 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_25_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf4), .Y(_20543_) );
	AOI21X1 AOI21X1_3140 ( .gnd(gnd), .vdd(vdd), .A(_20542_), .B(_20492__bF_buf4), .C(_20543_), .Y(_17349__25_) );
	INVX1 INVX1_3132 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_26_), .Y(_20544_) );
	OAI21X1 OAI21X1_4656 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_26_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf3), .Y(_20545_) );
	AOI21X1 AOI21X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_20544_), .B(_20492__bF_buf2), .C(_20545_), .Y(_17349__26_) );
	INVX1 INVX1_3133 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_27_), .Y(_20546_) );
	OAI21X1 OAI21X1_4657 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_27_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf2), .Y(_20547_) );
	AOI21X1 AOI21X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_20546_), .B(_20492__bF_buf0), .C(_20547_), .Y(_17349__27_) );
	INVX1 INVX1_3134 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_28_), .Y(_20548_) );
	OAI21X1 OAI21X1_4658 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_28_bF_buf4), .B(_20492__bF_buf7), .C(_19153__bF_buf1), .Y(_20549_) );
	AOI21X1 AOI21X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_20548_), .B(_20492__bF_buf6), .C(_20549_), .Y(_17349__28_) );
	INVX1 INVX1_3135 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_29_), .Y(_20550_) );
	OAI21X1 OAI21X1_4659 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_29_bF_buf4), .B(_20492__bF_buf5), .C(_19153__bF_buf0), .Y(_20551_) );
	AOI21X1 AOI21X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_20550_), .B(_20492__bF_buf4), .C(_20551_), .Y(_17349__29_) );
	INVX1 INVX1_3136 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_30_), .Y(_20552_) );
	OAI21X1 OAI21X1_4660 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_30_bF_buf4), .B(_20492__bF_buf3), .C(_19153__bF_buf98), .Y(_20553_) );
	AOI21X1 AOI21X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_20552_), .B(_20492__bF_buf2), .C(_20553_), .Y(_17349__30_) );
	INVX1 INVX1_3137 ( .gnd(gnd), .vdd(vdd), .A(registers_r1_31_), .Y(_20554_) );
	OAI21X1 OAI21X1_4661 ( .gnd(gnd), .vdd(vdd), .A(reg_dataIn_31_bF_buf4), .B(_20492__bF_buf1), .C(_19153__bF_buf97), .Y(_20555_) );
	AOI21X1 AOI21X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_20554_), .B(_20492__bF_buf0), .C(_20555_), .Y(_17349__31_) );
	INVX1 INVX1_3138 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_2_), .Y(_20556_) );
	NOR3X1 NOR3X1_203 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf5), .B(bLoc_frameOut_3_), .C(_20556_), .Y(_20557_) );
	INVX1 INVX1_3139 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .Y(_20558_) );
	NOR2X1 NOR2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_0_), .B(_20558_), .Y(_20559_) );
	NAND3X1 NAND3X1_3738 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_0_), .B(_20559__bF_buf5), .C(_20557__bF_buf7), .Y(_20560_) );
	NAND2X1 NAND2X1_3574 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .B(bLoc_frameOut_0_), .Y(_20561_) );
	INVX8 INVX8_74 ( .gnd(gnd), .vdd(vdd), .A(_20561_), .Y(_20562_) );
	NAND3X1 NAND3X1_3739 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_0_), .B(_20562__bF_buf5), .C(_20557__bF_buf6), .Y(_20563_) );
	NAND2X1 NAND2X1_3575 ( .gnd(gnd), .vdd(vdd), .A(_20560_), .B(_20563_), .Y(_20564_) );
	INVX4 INVX4_26 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf4), .Y(_20565_) );
	NOR2X1 NOR2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_3_), .B(bLoc_frameOut_2_), .Y(_20566_) );
	NAND3X1 NAND3X1_3740 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20566_), .C(_20559__bF_buf4), .Y(_20567_) );
	NAND3X1 NAND3X1_3741 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20566_), .C(_20562__bF_buf4), .Y(_20568_) );
	OAI22X1 OAI22X1_408 ( .gnd(gnd), .vdd(vdd), .A(_17379_), .B(_20568__bF_buf4), .C(_17380_), .D(_20567__bF_buf4), .Y(_20569_) );
	NOR2X1 NOR2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_20564_), .B(_20569_), .Y(_20570_) );
	INVX1 INVX1_3140 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_0_), .Y(_20571_) );
	NOR2X1 NOR2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .B(_20571_), .Y(_20572_) );
	INVX1 INVX1_3141 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_3_), .Y(_20573_) );
	NOR2X1 NOR2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_2_), .B(_20573_), .Y(_20574_) );
	NAND3X1 NAND3X1_3742 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20572_), .C(_20574__bF_buf7), .Y(_20575_) );
	NAND3X1 NAND3X1_3743 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20562__bF_buf3), .C(_20574__bF_buf6), .Y(_20576_) );
	OAI22X1 OAI22X1_409 ( .gnd(gnd), .vdd(vdd), .A(_17387_), .B(_20576__bF_buf4), .C(_17388_), .D(_20575__bF_buf4), .Y(_20577_) );
	NAND2X1 NAND2X1_3576 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_3_), .B(bLoc_frameOut_2_), .Y(_20578_) );
	INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(_20578_), .Y(_20579_) );
	NAND3X1 NAND3X1_3744 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20579_), .C(_20572_), .Y(_20580_) );
	NAND3X1 NAND3X1_3745 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20579_), .C(_20559__bF_buf3), .Y(_20581_) );
	OAI22X1 OAI22X1_410 ( .gnd(gnd), .vdd(vdd), .A(_17396_), .B(_20581__bF_buf4), .C(_17397_), .D(_20580__bF_buf4), .Y(_20582_) );
	NOR2X1 NOR2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_20582_), .B(_20577_), .Y(_20583_) );
	NAND2X1 NAND2X1_3577 ( .gnd(gnd), .vdd(vdd), .A(_20570_), .B(_20583_), .Y(_20584_) );
	NAND3X1 NAND3X1_3746 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf3), .B(_20566_), .C(_20559__bF_buf2), .Y(_20585_) );
	NAND3X1 NAND3X1_3747 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf2), .B(_20566_), .C(_20562__bF_buf2), .Y(_20586_) );
	OAI22X1 OAI22X1_411 ( .gnd(gnd), .vdd(vdd), .A(_17406_), .B(_20586__bF_buf4), .C(_17405_), .D(_20585__bF_buf4), .Y(_20587_) );
	NOR2X1 NOR2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_3_), .B(_20556_), .Y(_20588_) );
	NAND3X1 NAND3X1_3748 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf1), .B(_20572_), .C(_20588__bF_buf5), .Y(_20589_) );
	NOR3X1 NOR3X1_204 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .B(bLoc_frameOut_0_), .C(_20565_), .Y(_20590_) );
	NAND3X1 NAND3X1_3749 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_0_), .B(_20588__bF_buf4), .C(_20590__bF_buf7), .Y(_20591_) );
	OAI21X1 OAI21X1_4662 ( .gnd(gnd), .vdd(vdd), .A(_17410_), .B(_20589__bF_buf4), .C(_20591_), .Y(_20592_) );
	NOR2X1 NOR2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_20587_), .B(_20592_), .Y(_20593_) );
	NAND3X1 NAND3X1_3750 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf0), .B(_20579_), .C(_20559__bF_buf1), .Y(_20594_) );
	NOR2X1 NOR2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_20578_), .B(_20561_), .Y(_20595_) );
	NAND3X1 NAND3X1_3751 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_0_), .B(bLoc_frameOut_4_bF_buf6), .C(_20595__bF_buf4), .Y(_20596_) );
	OAI21X1 OAI21X1_4663 ( .gnd(gnd), .vdd(vdd), .A(_17417_), .B(_20594__bF_buf4), .C(_20596_), .Y(_20597_) );
	NAND3X1 NAND3X1_3752 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf5), .B(_20572_), .C(_20574__bF_buf5), .Y(_20598_) );
	NAND3X1 NAND3X1_3753 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_0_), .B(_20574__bF_buf4), .C(_20590__bF_buf6), .Y(_20599_) );
	OAI21X1 OAI21X1_4664 ( .gnd(gnd), .vdd(vdd), .A(_17422_), .B(_20598__bF_buf4), .C(_20599_), .Y(_20600_) );
	NOR2X1 NOR2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_20597_), .B(_20600_), .Y(_20601_) );
	NAND2X1 NAND2X1_3578 ( .gnd(gnd), .vdd(vdd), .A(_20601_), .B(_20593_), .Y(_20602_) );
	NOR2X1 NOR2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_20602_), .B(_20584_), .Y(_20603_) );
	NAND2X1 NAND2X1_3579 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_0_), .B(_20558_), .Y(_20604_) );
	INVX1 INVX1_3142 ( .gnd(gnd), .vdd(vdd), .A(_20566_), .Y(_20605_) );
	NOR3X1 NOR3X1_205 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf4), .B(_20604_), .C(_20605_), .Y(_20606_) );
	NOR3X1 NOR3X1_206 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf3), .B(bLoc_frameOut_1_), .C(bLoc_frameOut_0_), .Y(_20607_) );
	AND2X2 AND2X2_422 ( .gnd(gnd), .vdd(vdd), .A(_20607__bF_buf4), .B(_20579_), .Y(_20608_) );
	AOI22X1 AOI22X1_442 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_0_), .C(registers_r1_0_), .D(_20606__bF_buf4), .Y(_20609_) );
	AND2X2 AND2X2_423 ( .gnd(gnd), .vdd(vdd), .A(_20588__bF_buf3), .B(_20607__bF_buf3), .Y(_20610_) );
	AND2X2 AND2X2_424 ( .gnd(gnd), .vdd(vdd), .A(_20557__bF_buf5), .B(_20572_), .Y(_20611_) );
	AOI22X1 AOI22X1_443 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_0_), .C(registers_r5_0_), .D(_20611__bF_buf4), .Y(_20612_) );
	NAND2X1 NAND2X1_3580 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .B(_20571_), .Y(_20613_) );
	NAND2X1 NAND2X1_3581 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_3_), .B(_20556_), .Y(_20614_) );
	NOR3X1 NOR3X1_207 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf2), .B(_20613_), .C(_20614_), .Y(_20615_) );
	NAND3X1 NAND3X1_3754 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_0_), .B(_20607__bF_buf2), .C(_20574__bF_buf3), .Y(_20616_) );
	NAND3X1 NAND3X1_3755 ( .gnd(gnd), .vdd(vdd), .A(_20565_), .B(_20579_), .C(_20562__bF_buf1), .Y(_20617_) );
	OAI21X1 OAI21X1_4665 ( .gnd(gnd), .vdd(vdd), .A(_17441_), .B(_20617__bF_buf4), .C(_20616_), .Y(_20618_) );
	AOI21X1 AOI21X1_3147 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_0_), .B(_20615__bF_buf4), .C(_20618_), .Y(_20619_) );
	NAND3X1 NAND3X1_3756 ( .gnd(gnd), .vdd(vdd), .A(_20609_), .B(_20612_), .C(_20619_), .Y(_20620_) );
	NAND3X1 NAND3X1_3757 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf1), .B(_20588__bF_buf2), .C(_20559__bF_buf0), .Y(_20621_) );
	NAND3X1 NAND3X1_3758 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf0), .B(_20562__bF_buf0), .C(_20588__bF_buf1), .Y(_20622_) );
	OAI22X1 OAI22X1_412 ( .gnd(gnd), .vdd(vdd), .A(_17448_), .B(_20622__bF_buf4), .C(_17447_), .D(_20621__bF_buf4), .Y(_20623_) );
	NAND3X1 NAND3X1_3759 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf6), .B(_20566_), .C(_20572_), .Y(_20624_) );
	NOR2X1 NOR2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_1_), .B(bLoc_frameOut_0_), .Y(_20625_) );
	NAND3X1 NAND3X1_3760 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf5), .B(_20566_), .C(_20625_), .Y(_20626_) );
	OAI22X1 OAI22X1_413 ( .gnd(gnd), .vdd(vdd), .A(_17452_), .B(_20626__bF_buf4), .C(_17453_), .D(_20624__bF_buf4), .Y(_20627_) );
	NOR2X1 NOR2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_20627_), .B(_20623_), .Y(_20628_) );
	NAND3X1 NAND3X1_3761 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf4), .B(_20625_), .C(_20579_), .Y(_20629_) );
	NAND3X1 NAND3X1_3762 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf3), .B(_20579_), .C(_20572_), .Y(_20630_) );
	OAI22X1 OAI22X1_414 ( .gnd(gnd), .vdd(vdd), .A(_17459_), .B(_20629__bF_buf4), .C(_17460_), .D(_20630__bF_buf4), .Y(_20631_) );
	NAND3X1 NAND3X1_3763 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf2), .B(_20559__bF_buf5), .C(_20574__bF_buf2), .Y(_20632_) );
	NAND3X1 NAND3X1_3764 ( .gnd(gnd), .vdd(vdd), .A(bLoc_frameOut_4_bF_buf1), .B(_20562__bF_buf5), .C(_20574__bF_buf1), .Y(_20633_) );
	OAI22X1 OAI22X1_415 ( .gnd(gnd), .vdd(vdd), .A(_17465_), .B(_20633__bF_buf4), .C(_17464_), .D(_20632__bF_buf4), .Y(_20634_) );
	NOR2X1 NOR2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_20631_), .B(_20634_), .Y(_20635_) );
	NAND2X1 NAND2X1_3582 ( .gnd(gnd), .vdd(vdd), .A(_20628_), .B(_20635_), .Y(_20636_) );
	NOR2X1 NOR2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_20620_), .B(_20636_), .Y(_20637_) );
	NAND2X1 NAND2X1_3583 ( .gnd(gnd), .vdd(vdd), .A(_20637_), .B(_20603_), .Y(readB_regOut_0_) );
	NAND3X1 NAND3X1_3765 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_1_), .B(_20559__bF_buf4), .C(_20557__bF_buf4), .Y(_20638_) );
	NAND3X1 NAND3X1_3766 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_1_), .B(_20562__bF_buf4), .C(_20557__bF_buf3), .Y(_20639_) );
	NAND2X1 NAND2X1_3584 ( .gnd(gnd), .vdd(vdd), .A(_20638_), .B(_20639_), .Y(_20640_) );
	OAI22X1 OAI22X1_416 ( .gnd(gnd), .vdd(vdd), .A(_17475_), .B(_20568__bF_buf3), .C(_17476_), .D(_20567__bF_buf3), .Y(_20641_) );
	NOR2X1 NOR2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_20640_), .B(_20641_), .Y(_20642_) );
	OAI22X1 OAI22X1_417 ( .gnd(gnd), .vdd(vdd), .A(_17479_), .B(_20576__bF_buf3), .C(_17480_), .D(_20575__bF_buf3), .Y(_20643_) );
	OAI22X1 OAI22X1_418 ( .gnd(gnd), .vdd(vdd), .A(_17482_), .B(_20581__bF_buf3), .C(_17483_), .D(_20580__bF_buf3), .Y(_20644_) );
	NOR2X1 NOR2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_20644_), .B(_20643_), .Y(_20645_) );
	NAND2X1 NAND2X1_3585 ( .gnd(gnd), .vdd(vdd), .A(_20642_), .B(_20645_), .Y(_20646_) );
	OAI22X1 OAI22X1_419 ( .gnd(gnd), .vdd(vdd), .A(_17488_), .B(_20586__bF_buf3), .C(_17487_), .D(_20585__bF_buf3), .Y(_20647_) );
	NAND3X1 NAND3X1_3767 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_1_), .B(_20588__bF_buf0), .C(_20590__bF_buf5), .Y(_20648_) );
	OAI21X1 OAI21X1_4666 ( .gnd(gnd), .vdd(vdd), .A(_17490_), .B(_20589__bF_buf3), .C(_20648_), .Y(_20649_) );
	NOR2X1 NOR2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_20647_), .B(_20649_), .Y(_20650_) );
	NAND3X1 NAND3X1_3768 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_1_), .B(bLoc_frameOut_4_bF_buf0), .C(_20595__bF_buf3), .Y(_20651_) );
	OAI21X1 OAI21X1_4667 ( .gnd(gnd), .vdd(vdd), .A(_17494_), .B(_20594__bF_buf3), .C(_20651_), .Y(_20652_) );
	NAND3X1 NAND3X1_3769 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_1_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_20653_) );
	OAI21X1 OAI21X1_4668 ( .gnd(gnd), .vdd(vdd), .A(_17497_), .B(_20598__bF_buf3), .C(_20653_), .Y(_20654_) );
	NOR2X1 NOR2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_20652_), .B(_20654_), .Y(_20655_) );
	NAND2X1 NAND2X1_3586 ( .gnd(gnd), .vdd(vdd), .A(_20655_), .B(_20650_), .Y(_20656_) );
	NOR2X1 NOR2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_20656_), .B(_20646_), .Y(_20657_) );
	AOI22X1 AOI22X1_444 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_1_), .C(registers_r1_1_), .D(_20606__bF_buf3), .Y(_20658_) );
	AOI22X1 AOI22X1_445 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_1_), .C(registers_r5_1_), .D(_20611__bF_buf3), .Y(_20659_) );
	NAND3X1 NAND3X1_3770 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_1_), .B(_20607__bF_buf1), .C(_20574__bF_buf7), .Y(_20660_) );
	OAI21X1 OAI21X1_4669 ( .gnd(gnd), .vdd(vdd), .A(_17505_), .B(_20617__bF_buf3), .C(_20660_), .Y(_20661_) );
	AOI21X1 AOI21X1_3148 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_1_), .B(_20615__bF_buf3), .C(_20661_), .Y(_20662_) );
	NAND3X1 NAND3X1_3771 ( .gnd(gnd), .vdd(vdd), .A(_20658_), .B(_20659_), .C(_20662_), .Y(_20663_) );
	OAI22X1 OAI22X1_420 ( .gnd(gnd), .vdd(vdd), .A(_17511_), .B(_20622__bF_buf3), .C(_17510_), .D(_20621__bF_buf3), .Y(_20664_) );
	OAI22X1 OAI22X1_421 ( .gnd(gnd), .vdd(vdd), .A(_17513_), .B(_20626__bF_buf3), .C(_17514_), .D(_20624__bF_buf3), .Y(_20665_) );
	NOR2X1 NOR2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_20665_), .B(_20664_), .Y(_20666_) );
	OAI22X1 OAI22X1_422 ( .gnd(gnd), .vdd(vdd), .A(_17517_), .B(_20629__bF_buf3), .C(_17518_), .D(_20630__bF_buf3), .Y(_20667_) );
	OAI22X1 OAI22X1_423 ( .gnd(gnd), .vdd(vdd), .A(_17521_), .B(_20633__bF_buf3), .C(_17520_), .D(_20632__bF_buf3), .Y(_20668_) );
	NOR2X1 NOR2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_20667_), .B(_20668_), .Y(_20669_) );
	NAND2X1 NAND2X1_3587 ( .gnd(gnd), .vdd(vdd), .A(_20666_), .B(_20669_), .Y(_20670_) );
	NOR2X1 NOR2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_20663_), .B(_20670_), .Y(_20671_) );
	NAND2X1 NAND2X1_3588 ( .gnd(gnd), .vdd(vdd), .A(_20671_), .B(_20657_), .Y(readB_regOut_1_) );
	NAND3X1 NAND3X1_3772 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_2_), .B(_20559__bF_buf3), .C(_20557__bF_buf2), .Y(_20672_) );
	NAND3X1 NAND3X1_3773 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_2_), .B(_20562__bF_buf3), .C(_20557__bF_buf1), .Y(_20673_) );
	NAND2X1 NAND2X1_3589 ( .gnd(gnd), .vdd(vdd), .A(_20672_), .B(_20673_), .Y(_20674_) );
	OAI22X1 OAI22X1_424 ( .gnd(gnd), .vdd(vdd), .A(_17529_), .B(_20568__bF_buf2), .C(_17530_), .D(_20567__bF_buf2), .Y(_20675_) );
	NOR2X1 NOR2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_20674_), .B(_20675_), .Y(_20676_) );
	OAI22X1 OAI22X1_425 ( .gnd(gnd), .vdd(vdd), .A(_17533_), .B(_20576__bF_buf2), .C(_17534_), .D(_20575__bF_buf2), .Y(_20677_) );
	OAI22X1 OAI22X1_426 ( .gnd(gnd), .vdd(vdd), .A(_17536_), .B(_20581__bF_buf2), .C(_17537_), .D(_20580__bF_buf2), .Y(_20678_) );
	NOR2X1 NOR2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_20678_), .B(_20677_), .Y(_20679_) );
	NAND2X1 NAND2X1_3590 ( .gnd(gnd), .vdd(vdd), .A(_20676_), .B(_20679_), .Y(_20680_) );
	OAI22X1 OAI22X1_427 ( .gnd(gnd), .vdd(vdd), .A(_17542_), .B(_20586__bF_buf2), .C(_17541_), .D(_20585__bF_buf2), .Y(_20681_) );
	NAND3X1 NAND3X1_3774 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_2_), .B(_20588__bF_buf5), .C(_20590__bF_buf3), .Y(_20682_) );
	OAI21X1 OAI21X1_4670 ( .gnd(gnd), .vdd(vdd), .A(_17544_), .B(_20589__bF_buf2), .C(_20682_), .Y(_20683_) );
	NOR2X1 NOR2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_20681_), .B(_20683_), .Y(_20684_) );
	NAND3X1 NAND3X1_3775 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_2_), .B(bLoc_frameOut_4_bF_buf6), .C(_20595__bF_buf2), .Y(_20685_) );
	OAI21X1 OAI21X1_4671 ( .gnd(gnd), .vdd(vdd), .A(_17548_), .B(_20594__bF_buf2), .C(_20685_), .Y(_20686_) );
	NAND3X1 NAND3X1_3776 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_2_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_20687_) );
	OAI21X1 OAI21X1_4672 ( .gnd(gnd), .vdd(vdd), .A(_17551_), .B(_20598__bF_buf2), .C(_20687_), .Y(_20688_) );
	NOR2X1 NOR2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_20686_), .B(_20688_), .Y(_20689_) );
	NAND2X1 NAND2X1_3591 ( .gnd(gnd), .vdd(vdd), .A(_20689_), .B(_20684_), .Y(_20690_) );
	NOR2X1 NOR2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_20690_), .B(_20680_), .Y(_20691_) );
	AOI22X1 AOI22X1_446 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf2), .B(registers_a2_2_), .C(registers_r1_2_), .D(_20606__bF_buf2), .Y(_20692_) );
	AOI22X1 AOI22X1_447 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf2), .B(registers_r4_2_), .C(registers_r5_2_), .D(_20611__bF_buf2), .Y(_20693_) );
	NAND3X1 NAND3X1_3777 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_2_), .B(_20607__bF_buf0), .C(_20574__bF_buf5), .Y(_20694_) );
	OAI21X1 OAI21X1_4673 ( .gnd(gnd), .vdd(vdd), .A(_17559_), .B(_20617__bF_buf2), .C(_20694_), .Y(_20695_) );
	AOI21X1 AOI21X1_3149 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_2_), .B(_20615__bF_buf2), .C(_20695_), .Y(_20696_) );
	NAND3X1 NAND3X1_3778 ( .gnd(gnd), .vdd(vdd), .A(_20692_), .B(_20693_), .C(_20696_), .Y(_20697_) );
	OAI22X1 OAI22X1_428 ( .gnd(gnd), .vdd(vdd), .A(_17565_), .B(_20622__bF_buf2), .C(_17564_), .D(_20621__bF_buf2), .Y(_20698_) );
	OAI22X1 OAI22X1_429 ( .gnd(gnd), .vdd(vdd), .A(_17567_), .B(_20626__bF_buf2), .C(_17568_), .D(_20624__bF_buf2), .Y(_20699_) );
	NOR2X1 NOR2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_20699_), .B(_20698_), .Y(_20700_) );
	OAI22X1 OAI22X1_430 ( .gnd(gnd), .vdd(vdd), .A(_17571_), .B(_20629__bF_buf2), .C(_17572_), .D(_20630__bF_buf2), .Y(_20701_) );
	OAI22X1 OAI22X1_431 ( .gnd(gnd), .vdd(vdd), .A(_17575_), .B(_20633__bF_buf2), .C(_17574_), .D(_20632__bF_buf2), .Y(_20702_) );
	NOR2X1 NOR2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_20701_), .B(_20702_), .Y(_20703_) );
	NAND2X1 NAND2X1_3592 ( .gnd(gnd), .vdd(vdd), .A(_20700_), .B(_20703_), .Y(_20704_) );
	NOR2X1 NOR2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_20697_), .B(_20704_), .Y(_20705_) );
	NAND2X1 NAND2X1_3593 ( .gnd(gnd), .vdd(vdd), .A(_20705_), .B(_20691_), .Y(readB_regOut_2_) );
	NAND3X1 NAND3X1_3779 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_3_), .B(_20559__bF_buf2), .C(_20557__bF_buf0), .Y(_20706_) );
	NAND3X1 NAND3X1_3780 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_3_), .B(_20562__bF_buf2), .C(_20557__bF_buf7), .Y(_20707_) );
	NAND2X1 NAND2X1_3594 ( .gnd(gnd), .vdd(vdd), .A(_20706_), .B(_20707_), .Y(_20708_) );
	OAI22X1 OAI22X1_432 ( .gnd(gnd), .vdd(vdd), .A(_17583_), .B(_20568__bF_buf1), .C(_17584_), .D(_20567__bF_buf1), .Y(_20709_) );
	NOR2X1 NOR2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_20708_), .B(_20709_), .Y(_20710_) );
	OAI22X1 OAI22X1_433 ( .gnd(gnd), .vdd(vdd), .A(_17587_), .B(_20576__bF_buf1), .C(_17588_), .D(_20575__bF_buf1), .Y(_20711_) );
	OAI22X1 OAI22X1_434 ( .gnd(gnd), .vdd(vdd), .A(_17590_), .B(_20581__bF_buf1), .C(_17591_), .D(_20580__bF_buf1), .Y(_20712_) );
	NOR2X1 NOR2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_20712_), .B(_20711_), .Y(_20713_) );
	NAND2X1 NAND2X1_3595 ( .gnd(gnd), .vdd(vdd), .A(_20710_), .B(_20713_), .Y(_20714_) );
	OAI22X1 OAI22X1_435 ( .gnd(gnd), .vdd(vdd), .A(_17596_), .B(_20586__bF_buf1), .C(_17595_), .D(_20585__bF_buf1), .Y(_20715_) );
	NAND3X1 NAND3X1_3781 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_3_), .B(_20588__bF_buf4), .C(_20590__bF_buf1), .Y(_20716_) );
	OAI21X1 OAI21X1_4674 ( .gnd(gnd), .vdd(vdd), .A(_17598_), .B(_20589__bF_buf1), .C(_20716_), .Y(_20717_) );
	NOR2X1 NOR2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_20715_), .B(_20717_), .Y(_20718_) );
	NAND3X1 NAND3X1_3782 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_3_), .B(bLoc_frameOut_4_bF_buf5), .C(_20595__bF_buf1), .Y(_20719_) );
	OAI21X1 OAI21X1_4675 ( .gnd(gnd), .vdd(vdd), .A(_17602_), .B(_20594__bF_buf1), .C(_20719_), .Y(_20720_) );
	NAND3X1 NAND3X1_3783 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_3_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_20721_) );
	OAI21X1 OAI21X1_4676 ( .gnd(gnd), .vdd(vdd), .A(_17605_), .B(_20598__bF_buf1), .C(_20721_), .Y(_20722_) );
	NOR2X1 NOR2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_20720_), .B(_20722_), .Y(_20723_) );
	NAND2X1 NAND2X1_3596 ( .gnd(gnd), .vdd(vdd), .A(_20723_), .B(_20718_), .Y(_20724_) );
	NOR2X1 NOR2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_20724_), .B(_20714_), .Y(_20725_) );
	AOI22X1 AOI22X1_448 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf1), .B(registers_a2_3_), .C(registers_r1_3_), .D(_20606__bF_buf1), .Y(_20726_) );
	AOI22X1 AOI22X1_449 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf1), .B(registers_r4_3_), .C(registers_r5_3_), .D(_20611__bF_buf1), .Y(_20727_) );
	NAND3X1 NAND3X1_3784 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_3_), .B(_20607__bF_buf4), .C(_20574__bF_buf3), .Y(_20728_) );
	OAI21X1 OAI21X1_4677 ( .gnd(gnd), .vdd(vdd), .A(_17613_), .B(_20617__bF_buf1), .C(_20728_), .Y(_20729_) );
	AOI21X1 AOI21X1_3150 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_3_), .B(_20615__bF_buf1), .C(_20729_), .Y(_20730_) );
	NAND3X1 NAND3X1_3785 ( .gnd(gnd), .vdd(vdd), .A(_20726_), .B(_20727_), .C(_20730_), .Y(_20731_) );
	OAI22X1 OAI22X1_436 ( .gnd(gnd), .vdd(vdd), .A(_17619_), .B(_20622__bF_buf1), .C(_17618_), .D(_20621__bF_buf1), .Y(_20732_) );
	OAI22X1 OAI22X1_437 ( .gnd(gnd), .vdd(vdd), .A(_17621_), .B(_20626__bF_buf1), .C(_17622_), .D(_20624__bF_buf1), .Y(_20733_) );
	NOR2X1 NOR2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_20733_), .B(_20732_), .Y(_20734_) );
	OAI22X1 OAI22X1_438 ( .gnd(gnd), .vdd(vdd), .A(_17625_), .B(_20629__bF_buf1), .C(_17626_), .D(_20630__bF_buf1), .Y(_20735_) );
	OAI22X1 OAI22X1_439 ( .gnd(gnd), .vdd(vdd), .A(_17629_), .B(_20633__bF_buf1), .C(_17628_), .D(_20632__bF_buf1), .Y(_20736_) );
	NOR2X1 NOR2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_20735_), .B(_20736_), .Y(_20737_) );
	NAND2X1 NAND2X1_3597 ( .gnd(gnd), .vdd(vdd), .A(_20734_), .B(_20737_), .Y(_20738_) );
	NOR2X1 NOR2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_20731_), .B(_20738_), .Y(_20739_) );
	NAND2X1 NAND2X1_3598 ( .gnd(gnd), .vdd(vdd), .A(_20739_), .B(_20725_), .Y(readB_regOut_3_) );
	NAND3X1 NAND3X1_3786 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_4_), .B(_20559__bF_buf1), .C(_20557__bF_buf6), .Y(_20740_) );
	NAND3X1 NAND3X1_3787 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_4_), .B(_20562__bF_buf1), .C(_20557__bF_buf5), .Y(_20741_) );
	NAND2X1 NAND2X1_3599 ( .gnd(gnd), .vdd(vdd), .A(_20740_), .B(_20741_), .Y(_20742_) );
	OAI22X1 OAI22X1_440 ( .gnd(gnd), .vdd(vdd), .A(_17637_), .B(_20568__bF_buf0), .C(_17638_), .D(_20567__bF_buf0), .Y(_20743_) );
	NOR2X1 NOR2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_20742_), .B(_20743_), .Y(_20744_) );
	OAI22X1 OAI22X1_441 ( .gnd(gnd), .vdd(vdd), .A(_17641_), .B(_20576__bF_buf0), .C(_17642_), .D(_20575__bF_buf0), .Y(_20745_) );
	OAI22X1 OAI22X1_442 ( .gnd(gnd), .vdd(vdd), .A(_17644_), .B(_20581__bF_buf0), .C(_17645_), .D(_20580__bF_buf0), .Y(_20746_) );
	NOR2X1 NOR2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_20746_), .B(_20745_), .Y(_20747_) );
	NAND2X1 NAND2X1_3600 ( .gnd(gnd), .vdd(vdd), .A(_20744_), .B(_20747_), .Y(_20748_) );
	OAI22X1 OAI22X1_443 ( .gnd(gnd), .vdd(vdd), .A(_17650_), .B(_20586__bF_buf0), .C(_17649_), .D(_20585__bF_buf0), .Y(_20749_) );
	NAND3X1 NAND3X1_3788 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_4_), .B(_20588__bF_buf3), .C(_20590__bF_buf7), .Y(_20750_) );
	OAI21X1 OAI21X1_4678 ( .gnd(gnd), .vdd(vdd), .A(_17652_), .B(_20589__bF_buf0), .C(_20750_), .Y(_20751_) );
	NOR2X1 NOR2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_20749_), .B(_20751_), .Y(_20752_) );
	NAND3X1 NAND3X1_3789 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_4_), .B(bLoc_frameOut_4_bF_buf4), .C(_20595__bF_buf0), .Y(_20753_) );
	OAI21X1 OAI21X1_4679 ( .gnd(gnd), .vdd(vdd), .A(_17656_), .B(_20594__bF_buf0), .C(_20753_), .Y(_20754_) );
	NAND3X1 NAND3X1_3790 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_4_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_20755_) );
	OAI21X1 OAI21X1_4680 ( .gnd(gnd), .vdd(vdd), .A(_17659_), .B(_20598__bF_buf0), .C(_20755_), .Y(_20756_) );
	NOR2X1 NOR2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_20754_), .B(_20756_), .Y(_20757_) );
	NAND2X1 NAND2X1_3601 ( .gnd(gnd), .vdd(vdd), .A(_20757_), .B(_20752_), .Y(_20758_) );
	NOR2X1 NOR2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_20758_), .B(_20748_), .Y(_20759_) );
	AOI22X1 AOI22X1_450 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf0), .B(registers_a2_4_), .C(registers_r1_4_), .D(_20606__bF_buf0), .Y(_20760_) );
	AOI22X1 AOI22X1_451 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf0), .B(registers_r4_4_), .C(registers_r5_4_), .D(_20611__bF_buf0), .Y(_20761_) );
	NAND3X1 NAND3X1_3791 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_4_), .B(_20607__bF_buf3), .C(_20574__bF_buf1), .Y(_20762_) );
	OAI21X1 OAI21X1_4681 ( .gnd(gnd), .vdd(vdd), .A(_17667_), .B(_20617__bF_buf0), .C(_20762_), .Y(_20763_) );
	AOI21X1 AOI21X1_3151 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_4_), .B(_20615__bF_buf0), .C(_20763_), .Y(_20764_) );
	NAND3X1 NAND3X1_3792 ( .gnd(gnd), .vdd(vdd), .A(_20760_), .B(_20761_), .C(_20764_), .Y(_20765_) );
	OAI22X1 OAI22X1_444 ( .gnd(gnd), .vdd(vdd), .A(_17673_), .B(_20622__bF_buf0), .C(_17672_), .D(_20621__bF_buf0), .Y(_20766_) );
	OAI22X1 OAI22X1_445 ( .gnd(gnd), .vdd(vdd), .A(_17675_), .B(_20626__bF_buf0), .C(_17676_), .D(_20624__bF_buf0), .Y(_20767_) );
	NOR2X1 NOR2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_20767_), .B(_20766_), .Y(_20768_) );
	OAI22X1 OAI22X1_446 ( .gnd(gnd), .vdd(vdd), .A(_17679_), .B(_20629__bF_buf0), .C(_17680_), .D(_20630__bF_buf0), .Y(_20769_) );
	OAI22X1 OAI22X1_447 ( .gnd(gnd), .vdd(vdd), .A(_17683_), .B(_20633__bF_buf0), .C(_17682_), .D(_20632__bF_buf0), .Y(_20770_) );
	NOR2X1 NOR2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_20769_), .B(_20770_), .Y(_20771_) );
	NAND2X1 NAND2X1_3602 ( .gnd(gnd), .vdd(vdd), .A(_20768_), .B(_20771_), .Y(_20772_) );
	NOR2X1 NOR2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_20765_), .B(_20772_), .Y(_20773_) );
	NAND2X1 NAND2X1_3603 ( .gnd(gnd), .vdd(vdd), .A(_20773_), .B(_20759_), .Y(readB_regOut_4_) );
	NAND3X1 NAND3X1_3793 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_5_), .B(_20559__bF_buf0), .C(_20557__bF_buf4), .Y(_20774_) );
	NAND3X1 NAND3X1_3794 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_5_), .B(_20562__bF_buf0), .C(_20557__bF_buf3), .Y(_20775_) );
	NAND2X1 NAND2X1_3604 ( .gnd(gnd), .vdd(vdd), .A(_20774_), .B(_20775_), .Y(_20776_) );
	OAI22X1 OAI22X1_448 ( .gnd(gnd), .vdd(vdd), .A(_17691_), .B(_20568__bF_buf4), .C(_17692_), .D(_20567__bF_buf4), .Y(_20777_) );
	NOR2X1 NOR2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_20776_), .B(_20777_), .Y(_20778_) );
	OAI22X1 OAI22X1_449 ( .gnd(gnd), .vdd(vdd), .A(_17695_), .B(_20576__bF_buf4), .C(_17696_), .D(_20575__bF_buf4), .Y(_20779_) );
	OAI22X1 OAI22X1_450 ( .gnd(gnd), .vdd(vdd), .A(_17698_), .B(_20581__bF_buf4), .C(_17699_), .D(_20580__bF_buf4), .Y(_20780_) );
	NOR2X1 NOR2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_20780_), .B(_20779_), .Y(_20781_) );
	NAND2X1 NAND2X1_3605 ( .gnd(gnd), .vdd(vdd), .A(_20778_), .B(_20781_), .Y(_20782_) );
	OAI22X1 OAI22X1_451 ( .gnd(gnd), .vdd(vdd), .A(_17704_), .B(_20586__bF_buf4), .C(_17703_), .D(_20585__bF_buf4), .Y(_20783_) );
	NAND3X1 NAND3X1_3795 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_5_), .B(_20588__bF_buf2), .C(_20590__bF_buf5), .Y(_20784_) );
	OAI21X1 OAI21X1_4682 ( .gnd(gnd), .vdd(vdd), .A(_17706_), .B(_20589__bF_buf4), .C(_20784_), .Y(_20785_) );
	NOR2X1 NOR2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_20783_), .B(_20785_), .Y(_20786_) );
	NAND3X1 NAND3X1_3796 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_5_), .B(bLoc_frameOut_4_bF_buf3), .C(_20595__bF_buf4), .Y(_20787_) );
	OAI21X1 OAI21X1_4683 ( .gnd(gnd), .vdd(vdd), .A(_17710_), .B(_20594__bF_buf4), .C(_20787_), .Y(_20788_) );
	NAND3X1 NAND3X1_3797 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_5_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_20789_) );
	OAI21X1 OAI21X1_4684 ( .gnd(gnd), .vdd(vdd), .A(_17713_), .B(_20598__bF_buf4), .C(_20789_), .Y(_20790_) );
	NOR2X1 NOR2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_20788_), .B(_20790_), .Y(_20791_) );
	NAND2X1 NAND2X1_3606 ( .gnd(gnd), .vdd(vdd), .A(_20791_), .B(_20786_), .Y(_20792_) );
	NOR2X1 NOR2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_20792_), .B(_20782_), .Y(_20793_) );
	AOI22X1 AOI22X1_452 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_5_), .C(registers_r1_5_), .D(_20606__bF_buf4), .Y(_20794_) );
	AOI22X1 AOI22X1_453 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_5_), .C(registers_r5_5_), .D(_20611__bF_buf4), .Y(_20795_) );
	NAND3X1 NAND3X1_3798 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_5_), .B(_20607__bF_buf2), .C(_20574__bF_buf7), .Y(_20796_) );
	OAI21X1 OAI21X1_4685 ( .gnd(gnd), .vdd(vdd), .A(_17721_), .B(_20617__bF_buf4), .C(_20796_), .Y(_20797_) );
	AOI21X1 AOI21X1_3152 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_5_), .B(_20615__bF_buf4), .C(_20797_), .Y(_20798_) );
	NAND3X1 NAND3X1_3799 ( .gnd(gnd), .vdd(vdd), .A(_20794_), .B(_20795_), .C(_20798_), .Y(_20799_) );
	OAI22X1 OAI22X1_452 ( .gnd(gnd), .vdd(vdd), .A(_17727_), .B(_20622__bF_buf4), .C(_17726_), .D(_20621__bF_buf4), .Y(_20800_) );
	OAI22X1 OAI22X1_453 ( .gnd(gnd), .vdd(vdd), .A(_17729_), .B(_20626__bF_buf4), .C(_17730_), .D(_20624__bF_buf4), .Y(_20801_) );
	NOR2X1 NOR2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_20801_), .B(_20800_), .Y(_20802_) );
	OAI22X1 OAI22X1_454 ( .gnd(gnd), .vdd(vdd), .A(_17733_), .B(_20629__bF_buf4), .C(_17734_), .D(_20630__bF_buf4), .Y(_20803_) );
	OAI22X1 OAI22X1_455 ( .gnd(gnd), .vdd(vdd), .A(_17737_), .B(_20633__bF_buf4), .C(_17736_), .D(_20632__bF_buf4), .Y(_20804_) );
	NOR2X1 NOR2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_20803_), .B(_20804_), .Y(_20805_) );
	NAND2X1 NAND2X1_3607 ( .gnd(gnd), .vdd(vdd), .A(_20802_), .B(_20805_), .Y(_20806_) );
	NOR2X1 NOR2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_20799_), .B(_20806_), .Y(_20807_) );
	NAND2X1 NAND2X1_3608 ( .gnd(gnd), .vdd(vdd), .A(_20807_), .B(_20793_), .Y(readB_regOut_5_) );
	NAND3X1 NAND3X1_3800 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_6_), .B(_20559__bF_buf5), .C(_20557__bF_buf2), .Y(_20808_) );
	NAND3X1 NAND3X1_3801 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_6_), .B(_20562__bF_buf5), .C(_20557__bF_buf1), .Y(_20809_) );
	NAND2X1 NAND2X1_3609 ( .gnd(gnd), .vdd(vdd), .A(_20808_), .B(_20809_), .Y(_20810_) );
	OAI22X1 OAI22X1_456 ( .gnd(gnd), .vdd(vdd), .A(_17745_), .B(_20568__bF_buf3), .C(_17746_), .D(_20567__bF_buf3), .Y(_20811_) );
	NOR2X1 NOR2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_20810_), .B(_20811_), .Y(_20812_) );
	OAI22X1 OAI22X1_457 ( .gnd(gnd), .vdd(vdd), .A(_17749_), .B(_20576__bF_buf3), .C(_17750_), .D(_20575__bF_buf3), .Y(_20813_) );
	OAI22X1 OAI22X1_458 ( .gnd(gnd), .vdd(vdd), .A(_17752_), .B(_20581__bF_buf3), .C(_17753_), .D(_20580__bF_buf3), .Y(_20814_) );
	NOR2X1 NOR2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_20814_), .B(_20813_), .Y(_20815_) );
	NAND2X1 NAND2X1_3610 ( .gnd(gnd), .vdd(vdd), .A(_20812_), .B(_20815_), .Y(_20816_) );
	OAI22X1 OAI22X1_459 ( .gnd(gnd), .vdd(vdd), .A(_17758_), .B(_20586__bF_buf3), .C(_17757_), .D(_20585__bF_buf3), .Y(_20817_) );
	NAND3X1 NAND3X1_3802 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_6_), .B(_20588__bF_buf1), .C(_20590__bF_buf3), .Y(_20818_) );
	OAI21X1 OAI21X1_4686 ( .gnd(gnd), .vdd(vdd), .A(_17760_), .B(_20589__bF_buf3), .C(_20818_), .Y(_20819_) );
	NOR2X1 NOR2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_20817_), .B(_20819_), .Y(_20820_) );
	NAND3X1 NAND3X1_3803 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_6_), .B(bLoc_frameOut_4_bF_buf2), .C(_20595__bF_buf3), .Y(_20821_) );
	OAI21X1 OAI21X1_4687 ( .gnd(gnd), .vdd(vdd), .A(_17764_), .B(_20594__bF_buf3), .C(_20821_), .Y(_20822_) );
	NAND3X1 NAND3X1_3804 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_6_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_20823_) );
	OAI21X1 OAI21X1_4688 ( .gnd(gnd), .vdd(vdd), .A(_17767_), .B(_20598__bF_buf3), .C(_20823_), .Y(_20824_) );
	NOR2X1 NOR2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_20822_), .B(_20824_), .Y(_20825_) );
	NAND2X1 NAND2X1_3611 ( .gnd(gnd), .vdd(vdd), .A(_20825_), .B(_20820_), .Y(_20826_) );
	NOR2X1 NOR2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_20826_), .B(_20816_), .Y(_20827_) );
	AOI22X1 AOI22X1_454 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_6_), .C(registers_r1_6_), .D(_20606__bF_buf3), .Y(_20828_) );
	AOI22X1 AOI22X1_455 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_6_), .C(registers_r5_6_), .D(_20611__bF_buf3), .Y(_20829_) );
	NAND3X1 NAND3X1_3805 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_6_), .B(_20607__bF_buf1), .C(_20574__bF_buf5), .Y(_20830_) );
	OAI21X1 OAI21X1_4689 ( .gnd(gnd), .vdd(vdd), .A(_17775_), .B(_20617__bF_buf3), .C(_20830_), .Y(_20831_) );
	AOI21X1 AOI21X1_3153 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_6_), .B(_20615__bF_buf3), .C(_20831_), .Y(_20832_) );
	NAND3X1 NAND3X1_3806 ( .gnd(gnd), .vdd(vdd), .A(_20828_), .B(_20829_), .C(_20832_), .Y(_20833_) );
	OAI22X1 OAI22X1_460 ( .gnd(gnd), .vdd(vdd), .A(_17781_), .B(_20622__bF_buf3), .C(_17780_), .D(_20621__bF_buf3), .Y(_20834_) );
	OAI22X1 OAI22X1_461 ( .gnd(gnd), .vdd(vdd), .A(_17783_), .B(_20626__bF_buf3), .C(_17784_), .D(_20624__bF_buf3), .Y(_20835_) );
	NOR2X1 NOR2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_20835_), .B(_20834_), .Y(_20836_) );
	OAI22X1 OAI22X1_462 ( .gnd(gnd), .vdd(vdd), .A(_17787_), .B(_20629__bF_buf3), .C(_17788_), .D(_20630__bF_buf3), .Y(_20837_) );
	OAI22X1 OAI22X1_463 ( .gnd(gnd), .vdd(vdd), .A(_17791_), .B(_20633__bF_buf3), .C(_17790_), .D(_20632__bF_buf3), .Y(_20838_) );
	NOR2X1 NOR2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_20837_), .B(_20838_), .Y(_20839_) );
	NAND2X1 NAND2X1_3612 ( .gnd(gnd), .vdd(vdd), .A(_20836_), .B(_20839_), .Y(_20840_) );
	NOR2X1 NOR2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_20833_), .B(_20840_), .Y(_20841_) );
	NAND2X1 NAND2X1_3613 ( .gnd(gnd), .vdd(vdd), .A(_20841_), .B(_20827_), .Y(readB_regOut_6_) );
	NAND3X1 NAND3X1_3807 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_7_), .B(_20559__bF_buf4), .C(_20557__bF_buf0), .Y(_20842_) );
	NAND3X1 NAND3X1_3808 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_7_), .B(_20562__bF_buf4), .C(_20557__bF_buf7), .Y(_20843_) );
	NAND2X1 NAND2X1_3614 ( .gnd(gnd), .vdd(vdd), .A(_20842_), .B(_20843_), .Y(_20844_) );
	OAI22X1 OAI22X1_464 ( .gnd(gnd), .vdd(vdd), .A(_17799_), .B(_20568__bF_buf2), .C(_17800_), .D(_20567__bF_buf2), .Y(_20845_) );
	NOR2X1 NOR2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_20844_), .B(_20845_), .Y(_20846_) );
	OAI22X1 OAI22X1_465 ( .gnd(gnd), .vdd(vdd), .A(_17803_), .B(_20576__bF_buf2), .C(_17804_), .D(_20575__bF_buf2), .Y(_20847_) );
	OAI22X1 OAI22X1_466 ( .gnd(gnd), .vdd(vdd), .A(_17806_), .B(_20581__bF_buf2), .C(_17807_), .D(_20580__bF_buf2), .Y(_20848_) );
	NOR2X1 NOR2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_20848_), .B(_20847_), .Y(_20849_) );
	NAND2X1 NAND2X1_3615 ( .gnd(gnd), .vdd(vdd), .A(_20846_), .B(_20849_), .Y(_20850_) );
	OAI22X1 OAI22X1_467 ( .gnd(gnd), .vdd(vdd), .A(_17812_), .B(_20586__bF_buf2), .C(_17811_), .D(_20585__bF_buf2), .Y(_20851_) );
	NAND3X1 NAND3X1_3809 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_7_), .B(_20588__bF_buf0), .C(_20590__bF_buf1), .Y(_20852_) );
	OAI21X1 OAI21X1_4690 ( .gnd(gnd), .vdd(vdd), .A(_17814_), .B(_20589__bF_buf2), .C(_20852_), .Y(_20853_) );
	NOR2X1 NOR2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_20851_), .B(_20853_), .Y(_20854_) );
	NAND3X1 NAND3X1_3810 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_7_), .B(bLoc_frameOut_4_bF_buf1), .C(_20595__bF_buf2), .Y(_20855_) );
	OAI21X1 OAI21X1_4691 ( .gnd(gnd), .vdd(vdd), .A(_17818_), .B(_20594__bF_buf2), .C(_20855_), .Y(_20856_) );
	NAND3X1 NAND3X1_3811 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_7_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_20857_) );
	OAI21X1 OAI21X1_4692 ( .gnd(gnd), .vdd(vdd), .A(_17821_), .B(_20598__bF_buf2), .C(_20857_), .Y(_20858_) );
	NOR2X1 NOR2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_20856_), .B(_20858_), .Y(_20859_) );
	NAND2X1 NAND2X1_3616 ( .gnd(gnd), .vdd(vdd), .A(_20859_), .B(_20854_), .Y(_20860_) );
	NOR2X1 NOR2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_20860_), .B(_20850_), .Y(_20861_) );
	AOI22X1 AOI22X1_456 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf2), .B(registers_a2_7_), .C(registers_r1_7_), .D(_20606__bF_buf2), .Y(_20862_) );
	AOI22X1 AOI22X1_457 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf2), .B(registers_r4_7_), .C(registers_r5_7_), .D(_20611__bF_buf2), .Y(_20863_) );
	NAND3X1 NAND3X1_3812 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_7_), .B(_20607__bF_buf0), .C(_20574__bF_buf3), .Y(_20864_) );
	OAI21X1 OAI21X1_4693 ( .gnd(gnd), .vdd(vdd), .A(_17829_), .B(_20617__bF_buf2), .C(_20864_), .Y(_20865_) );
	AOI21X1 AOI21X1_3154 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_7_), .B(_20615__bF_buf2), .C(_20865_), .Y(_20866_) );
	NAND3X1 NAND3X1_3813 ( .gnd(gnd), .vdd(vdd), .A(_20862_), .B(_20863_), .C(_20866_), .Y(_20867_) );
	OAI22X1 OAI22X1_468 ( .gnd(gnd), .vdd(vdd), .A(_17835_), .B(_20622__bF_buf2), .C(_17834_), .D(_20621__bF_buf2), .Y(_20868_) );
	OAI22X1 OAI22X1_469 ( .gnd(gnd), .vdd(vdd), .A(_17837_), .B(_20626__bF_buf2), .C(_17838_), .D(_20624__bF_buf2), .Y(_20869_) );
	NOR2X1 NOR2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_20869_), .B(_20868_), .Y(_20870_) );
	OAI22X1 OAI22X1_470 ( .gnd(gnd), .vdd(vdd), .A(_17841_), .B(_20629__bF_buf2), .C(_17842_), .D(_20630__bF_buf2), .Y(_20871_) );
	OAI22X1 OAI22X1_471 ( .gnd(gnd), .vdd(vdd), .A(_17845_), .B(_20633__bF_buf2), .C(_17844_), .D(_20632__bF_buf2), .Y(_20872_) );
	NOR2X1 NOR2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_20871_), .B(_20872_), .Y(_20873_) );
	NAND2X1 NAND2X1_3617 ( .gnd(gnd), .vdd(vdd), .A(_20870_), .B(_20873_), .Y(_20874_) );
	NOR2X1 NOR2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_20867_), .B(_20874_), .Y(_20875_) );
	NAND2X1 NAND2X1_3618 ( .gnd(gnd), .vdd(vdd), .A(_20875_), .B(_20861_), .Y(readB_regOut_7_) );
	NAND3X1 NAND3X1_3814 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_8_), .B(_20559__bF_buf3), .C(_20557__bF_buf6), .Y(_20876_) );
	NAND3X1 NAND3X1_3815 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_8_), .B(_20562__bF_buf3), .C(_20557__bF_buf5), .Y(_20877_) );
	NAND2X1 NAND2X1_3619 ( .gnd(gnd), .vdd(vdd), .A(_20876_), .B(_20877_), .Y(_20878_) );
	OAI22X1 OAI22X1_472 ( .gnd(gnd), .vdd(vdd), .A(_17853_), .B(_20568__bF_buf1), .C(_17854_), .D(_20567__bF_buf1), .Y(_20879_) );
	NOR2X1 NOR2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_20878_), .B(_20879_), .Y(_20880_) );
	OAI22X1 OAI22X1_473 ( .gnd(gnd), .vdd(vdd), .A(_17857_), .B(_20576__bF_buf1), .C(_17858_), .D(_20575__bF_buf1), .Y(_20881_) );
	OAI22X1 OAI22X1_474 ( .gnd(gnd), .vdd(vdd), .A(_17860_), .B(_20581__bF_buf1), .C(_17861_), .D(_20580__bF_buf1), .Y(_20882_) );
	NOR2X1 NOR2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_20882_), .B(_20881_), .Y(_20883_) );
	NAND2X1 NAND2X1_3620 ( .gnd(gnd), .vdd(vdd), .A(_20880_), .B(_20883_), .Y(_20884_) );
	OAI22X1 OAI22X1_475 ( .gnd(gnd), .vdd(vdd), .A(_17866_), .B(_20586__bF_buf1), .C(_17865_), .D(_20585__bF_buf1), .Y(_20885_) );
	NAND3X1 NAND3X1_3816 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_8_), .B(_20588__bF_buf5), .C(_20590__bF_buf7), .Y(_20886_) );
	OAI21X1 OAI21X1_4694 ( .gnd(gnd), .vdd(vdd), .A(_17868_), .B(_20589__bF_buf1), .C(_20886_), .Y(_20887_) );
	NOR2X1 NOR2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_20885_), .B(_20887_), .Y(_20888_) );
	NAND3X1 NAND3X1_3817 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_8_), .B(bLoc_frameOut_4_bF_buf0), .C(_20595__bF_buf1), .Y(_20889_) );
	OAI21X1 OAI21X1_4695 ( .gnd(gnd), .vdd(vdd), .A(_17872_), .B(_20594__bF_buf1), .C(_20889_), .Y(_20890_) );
	NAND3X1 NAND3X1_3818 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_8_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_20891_) );
	OAI21X1 OAI21X1_4696 ( .gnd(gnd), .vdd(vdd), .A(_17875_), .B(_20598__bF_buf1), .C(_20891_), .Y(_20892_) );
	NOR2X1 NOR2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_20890_), .B(_20892_), .Y(_20893_) );
	NAND2X1 NAND2X1_3621 ( .gnd(gnd), .vdd(vdd), .A(_20893_), .B(_20888_), .Y(_20894_) );
	NOR2X1 NOR2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_20894_), .B(_20884_), .Y(_20895_) );
	AOI22X1 AOI22X1_458 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf1), .B(registers_a2_8_), .C(registers_r1_8_), .D(_20606__bF_buf1), .Y(_20896_) );
	AOI22X1 AOI22X1_459 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf1), .B(registers_r4_8_), .C(registers_r5_8_), .D(_20611__bF_buf1), .Y(_20897_) );
	NAND3X1 NAND3X1_3819 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_8_), .B(_20607__bF_buf4), .C(_20574__bF_buf1), .Y(_20898_) );
	OAI21X1 OAI21X1_4697 ( .gnd(gnd), .vdd(vdd), .A(_17883_), .B(_20617__bF_buf1), .C(_20898_), .Y(_20899_) );
	AOI21X1 AOI21X1_3155 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_8_), .B(_20615__bF_buf1), .C(_20899_), .Y(_20900_) );
	NAND3X1 NAND3X1_3820 ( .gnd(gnd), .vdd(vdd), .A(_20896_), .B(_20897_), .C(_20900_), .Y(_20901_) );
	OAI22X1 OAI22X1_476 ( .gnd(gnd), .vdd(vdd), .A(_17889_), .B(_20622__bF_buf1), .C(_17888_), .D(_20621__bF_buf1), .Y(_20902_) );
	OAI22X1 OAI22X1_477 ( .gnd(gnd), .vdd(vdd), .A(_17891_), .B(_20626__bF_buf1), .C(_17892_), .D(_20624__bF_buf1), .Y(_20903_) );
	NOR2X1 NOR2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_20903_), .B(_20902_), .Y(_20904_) );
	OAI22X1 OAI22X1_478 ( .gnd(gnd), .vdd(vdd), .A(_17895_), .B(_20629__bF_buf1), .C(_17896_), .D(_20630__bF_buf1), .Y(_20905_) );
	OAI22X1 OAI22X1_479 ( .gnd(gnd), .vdd(vdd), .A(_17899_), .B(_20633__bF_buf1), .C(_17898_), .D(_20632__bF_buf1), .Y(_20906_) );
	NOR2X1 NOR2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_20905_), .B(_20906_), .Y(_20907_) );
	NAND2X1 NAND2X1_3622 ( .gnd(gnd), .vdd(vdd), .A(_20904_), .B(_20907_), .Y(_20908_) );
	NOR2X1 NOR2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_20901_), .B(_20908_), .Y(_20909_) );
	NAND2X1 NAND2X1_3623 ( .gnd(gnd), .vdd(vdd), .A(_20909_), .B(_20895_), .Y(readB_regOut_8_) );
	NAND3X1 NAND3X1_3821 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_9_), .B(_20559__bF_buf2), .C(_20557__bF_buf4), .Y(_20910_) );
	NAND3X1 NAND3X1_3822 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_9_), .B(_20562__bF_buf2), .C(_20557__bF_buf3), .Y(_20911_) );
	NAND2X1 NAND2X1_3624 ( .gnd(gnd), .vdd(vdd), .A(_20910_), .B(_20911_), .Y(_20912_) );
	OAI22X1 OAI22X1_480 ( .gnd(gnd), .vdd(vdd), .A(_17907_), .B(_20568__bF_buf0), .C(_17908_), .D(_20567__bF_buf0), .Y(_20913_) );
	NOR2X1 NOR2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_20912_), .B(_20913_), .Y(_20914_) );
	OAI22X1 OAI22X1_481 ( .gnd(gnd), .vdd(vdd), .A(_17911_), .B(_20576__bF_buf0), .C(_17912_), .D(_20575__bF_buf0), .Y(_20915_) );
	OAI22X1 OAI22X1_482 ( .gnd(gnd), .vdd(vdd), .A(_17914_), .B(_20581__bF_buf0), .C(_17915_), .D(_20580__bF_buf0), .Y(_20916_) );
	NOR2X1 NOR2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_20916_), .B(_20915_), .Y(_20917_) );
	NAND2X1 NAND2X1_3625 ( .gnd(gnd), .vdd(vdd), .A(_20914_), .B(_20917_), .Y(_20918_) );
	OAI22X1 OAI22X1_483 ( .gnd(gnd), .vdd(vdd), .A(_17920_), .B(_20586__bF_buf0), .C(_17919_), .D(_20585__bF_buf0), .Y(_20919_) );
	NAND3X1 NAND3X1_3823 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_9_), .B(_20588__bF_buf4), .C(_20590__bF_buf5), .Y(_20920_) );
	OAI21X1 OAI21X1_4698 ( .gnd(gnd), .vdd(vdd), .A(_17922_), .B(_20589__bF_buf0), .C(_20920_), .Y(_20921_) );
	NOR2X1 NOR2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_20919_), .B(_20921_), .Y(_20922_) );
	NAND3X1 NAND3X1_3824 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_9_), .B(bLoc_frameOut_4_bF_buf6), .C(_20595__bF_buf0), .Y(_20923_) );
	OAI21X1 OAI21X1_4699 ( .gnd(gnd), .vdd(vdd), .A(_17926_), .B(_20594__bF_buf0), .C(_20923_), .Y(_20924_) );
	NAND3X1 NAND3X1_3825 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_9_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_20925_) );
	OAI21X1 OAI21X1_4700 ( .gnd(gnd), .vdd(vdd), .A(_17929_), .B(_20598__bF_buf0), .C(_20925_), .Y(_20926_) );
	NOR2X1 NOR2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_20924_), .B(_20926_), .Y(_20927_) );
	NAND2X1 NAND2X1_3626 ( .gnd(gnd), .vdd(vdd), .A(_20927_), .B(_20922_), .Y(_20928_) );
	NOR2X1 NOR2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_20928_), .B(_20918_), .Y(_20929_) );
	AOI22X1 AOI22X1_460 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf0), .B(registers_a2_9_), .C(registers_r1_9_), .D(_20606__bF_buf0), .Y(_20930_) );
	AOI22X1 AOI22X1_461 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf0), .B(registers_r4_9_), .C(registers_r5_9_), .D(_20611__bF_buf0), .Y(_20931_) );
	NAND3X1 NAND3X1_3826 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_9_), .B(_20607__bF_buf3), .C(_20574__bF_buf7), .Y(_20932_) );
	OAI21X1 OAI21X1_4701 ( .gnd(gnd), .vdd(vdd), .A(_17937_), .B(_20617__bF_buf0), .C(_20932_), .Y(_20933_) );
	AOI21X1 AOI21X1_3156 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_9_), .B(_20615__bF_buf0), .C(_20933_), .Y(_20934_) );
	NAND3X1 NAND3X1_3827 ( .gnd(gnd), .vdd(vdd), .A(_20930_), .B(_20931_), .C(_20934_), .Y(_20935_) );
	OAI22X1 OAI22X1_484 ( .gnd(gnd), .vdd(vdd), .A(_17943_), .B(_20622__bF_buf0), .C(_17942_), .D(_20621__bF_buf0), .Y(_20936_) );
	OAI22X1 OAI22X1_485 ( .gnd(gnd), .vdd(vdd), .A(_17945_), .B(_20626__bF_buf0), .C(_17946_), .D(_20624__bF_buf0), .Y(_20937_) );
	NOR2X1 NOR2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_20937_), .B(_20936_), .Y(_20938_) );
	OAI22X1 OAI22X1_486 ( .gnd(gnd), .vdd(vdd), .A(_17949_), .B(_20629__bF_buf0), .C(_17950_), .D(_20630__bF_buf0), .Y(_20939_) );
	OAI22X1 OAI22X1_487 ( .gnd(gnd), .vdd(vdd), .A(_17953_), .B(_20633__bF_buf0), .C(_17952_), .D(_20632__bF_buf0), .Y(_20940_) );
	NOR2X1 NOR2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_20939_), .B(_20940_), .Y(_20941_) );
	NAND2X1 NAND2X1_3627 ( .gnd(gnd), .vdd(vdd), .A(_20938_), .B(_20941_), .Y(_20942_) );
	NOR2X1 NOR2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_20935_), .B(_20942_), .Y(_20943_) );
	NAND2X1 NAND2X1_3628 ( .gnd(gnd), .vdd(vdd), .A(_20943_), .B(_20929_), .Y(readB_regOut_9_) );
	NAND3X1 NAND3X1_3828 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_10_), .B(_20559__bF_buf1), .C(_20557__bF_buf2), .Y(_20944_) );
	NAND3X1 NAND3X1_3829 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_10_), .B(_20562__bF_buf1), .C(_20557__bF_buf1), .Y(_20945_) );
	NAND2X1 NAND2X1_3629 ( .gnd(gnd), .vdd(vdd), .A(_20944_), .B(_20945_), .Y(_20946_) );
	OAI22X1 OAI22X1_488 ( .gnd(gnd), .vdd(vdd), .A(_17961_), .B(_20568__bF_buf4), .C(_17962_), .D(_20567__bF_buf4), .Y(_20947_) );
	NOR2X1 NOR2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_20946_), .B(_20947_), .Y(_20948_) );
	OAI22X1 OAI22X1_489 ( .gnd(gnd), .vdd(vdd), .A(_17965_), .B(_20576__bF_buf4), .C(_17966_), .D(_20575__bF_buf4), .Y(_20949_) );
	OAI22X1 OAI22X1_490 ( .gnd(gnd), .vdd(vdd), .A(_17968_), .B(_20581__bF_buf4), .C(_17969_), .D(_20580__bF_buf4), .Y(_20950_) );
	NOR2X1 NOR2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_20950_), .B(_20949_), .Y(_20951_) );
	NAND2X1 NAND2X1_3630 ( .gnd(gnd), .vdd(vdd), .A(_20948_), .B(_20951_), .Y(_20952_) );
	OAI22X1 OAI22X1_491 ( .gnd(gnd), .vdd(vdd), .A(_17974_), .B(_20586__bF_buf4), .C(_17973_), .D(_20585__bF_buf4), .Y(_20953_) );
	NAND3X1 NAND3X1_3830 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_10_), .B(_20588__bF_buf3), .C(_20590__bF_buf3), .Y(_20954_) );
	OAI21X1 OAI21X1_4702 ( .gnd(gnd), .vdd(vdd), .A(_17976_), .B(_20589__bF_buf4), .C(_20954_), .Y(_20955_) );
	NOR2X1 NOR2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_20953_), .B(_20955_), .Y(_20956_) );
	NAND3X1 NAND3X1_3831 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_10_), .B(bLoc_frameOut_4_bF_buf5), .C(_20595__bF_buf4), .Y(_20957_) );
	OAI21X1 OAI21X1_4703 ( .gnd(gnd), .vdd(vdd), .A(_17980_), .B(_20594__bF_buf4), .C(_20957_), .Y(_20958_) );
	NAND3X1 NAND3X1_3832 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_10_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_20959_) );
	OAI21X1 OAI21X1_4704 ( .gnd(gnd), .vdd(vdd), .A(_17983_), .B(_20598__bF_buf4), .C(_20959_), .Y(_20960_) );
	NOR2X1 NOR2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_20958_), .B(_20960_), .Y(_20961_) );
	NAND2X1 NAND2X1_3631 ( .gnd(gnd), .vdd(vdd), .A(_20961_), .B(_20956_), .Y(_20962_) );
	NOR2X1 NOR2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_20962_), .B(_20952_), .Y(_20963_) );
	AOI22X1 AOI22X1_462 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_10_), .C(registers_r1_10_), .D(_20606__bF_buf4), .Y(_20964_) );
	AOI22X1 AOI22X1_463 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_10_), .C(registers_r5_10_), .D(_20611__bF_buf4), .Y(_20965_) );
	NAND3X1 NAND3X1_3833 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_10_), .B(_20607__bF_buf2), .C(_20574__bF_buf5), .Y(_20966_) );
	OAI21X1 OAI21X1_4705 ( .gnd(gnd), .vdd(vdd), .A(_17991_), .B(_20617__bF_buf4), .C(_20966_), .Y(_20967_) );
	AOI21X1 AOI21X1_3157 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_10_), .B(_20615__bF_buf4), .C(_20967_), .Y(_20968_) );
	NAND3X1 NAND3X1_3834 ( .gnd(gnd), .vdd(vdd), .A(_20964_), .B(_20965_), .C(_20968_), .Y(_20969_) );
	OAI22X1 OAI22X1_492 ( .gnd(gnd), .vdd(vdd), .A(_17997_), .B(_20622__bF_buf4), .C(_17996_), .D(_20621__bF_buf4), .Y(_20970_) );
	OAI22X1 OAI22X1_493 ( .gnd(gnd), .vdd(vdd), .A(_17999_), .B(_20626__bF_buf4), .C(_18000_), .D(_20624__bF_buf4), .Y(_20971_) );
	NOR2X1 NOR2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_20971_), .B(_20970_), .Y(_20972_) );
	OAI22X1 OAI22X1_494 ( .gnd(gnd), .vdd(vdd), .A(_18003_), .B(_20629__bF_buf4), .C(_18004_), .D(_20630__bF_buf4), .Y(_20973_) );
	OAI22X1 OAI22X1_495 ( .gnd(gnd), .vdd(vdd), .A(_18007_), .B(_20633__bF_buf4), .C(_18006_), .D(_20632__bF_buf4), .Y(_20974_) );
	NOR2X1 NOR2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_20973_), .B(_20974_), .Y(_20975_) );
	NAND2X1 NAND2X1_3632 ( .gnd(gnd), .vdd(vdd), .A(_20972_), .B(_20975_), .Y(_20976_) );
	NOR2X1 NOR2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_20969_), .B(_20976_), .Y(_20977_) );
	NAND2X1 NAND2X1_3633 ( .gnd(gnd), .vdd(vdd), .A(_20977_), .B(_20963_), .Y(readB_regOut_10_) );
	NAND3X1 NAND3X1_3835 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_11_), .B(_20559__bF_buf0), .C(_20557__bF_buf0), .Y(_20978_) );
	NAND3X1 NAND3X1_3836 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_11_), .B(_20562__bF_buf0), .C(_20557__bF_buf7), .Y(_20979_) );
	NAND2X1 NAND2X1_3634 ( .gnd(gnd), .vdd(vdd), .A(_20978_), .B(_20979_), .Y(_20980_) );
	OAI22X1 OAI22X1_496 ( .gnd(gnd), .vdd(vdd), .A(_18015_), .B(_20568__bF_buf3), .C(_18016_), .D(_20567__bF_buf3), .Y(_20981_) );
	NOR2X1 NOR2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_20980_), .B(_20981_), .Y(_20982_) );
	OAI22X1 OAI22X1_497 ( .gnd(gnd), .vdd(vdd), .A(_18019_), .B(_20576__bF_buf3), .C(_18020_), .D(_20575__bF_buf3), .Y(_20983_) );
	OAI22X1 OAI22X1_498 ( .gnd(gnd), .vdd(vdd), .A(_18022_), .B(_20581__bF_buf3), .C(_18023_), .D(_20580__bF_buf3), .Y(_20984_) );
	NOR2X1 NOR2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_20984_), .B(_20983_), .Y(_20985_) );
	NAND2X1 NAND2X1_3635 ( .gnd(gnd), .vdd(vdd), .A(_20982_), .B(_20985_), .Y(_20986_) );
	OAI22X1 OAI22X1_499 ( .gnd(gnd), .vdd(vdd), .A(_18028_), .B(_20586__bF_buf3), .C(_18027_), .D(_20585__bF_buf3), .Y(_20987_) );
	NAND3X1 NAND3X1_3837 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_11_), .B(_20588__bF_buf2), .C(_20590__bF_buf1), .Y(_20988_) );
	OAI21X1 OAI21X1_4706 ( .gnd(gnd), .vdd(vdd), .A(_18030_), .B(_20589__bF_buf3), .C(_20988_), .Y(_20989_) );
	NOR2X1 NOR2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_20987_), .B(_20989_), .Y(_20990_) );
	NAND3X1 NAND3X1_3838 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_11_), .B(bLoc_frameOut_4_bF_buf4), .C(_20595__bF_buf3), .Y(_20991_) );
	OAI21X1 OAI21X1_4707 ( .gnd(gnd), .vdd(vdd), .A(_18034_), .B(_20594__bF_buf3), .C(_20991_), .Y(_20992_) );
	NAND3X1 NAND3X1_3839 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_11_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_20993_) );
	OAI21X1 OAI21X1_4708 ( .gnd(gnd), .vdd(vdd), .A(_18037_), .B(_20598__bF_buf3), .C(_20993_), .Y(_20994_) );
	NOR2X1 NOR2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_20992_), .B(_20994_), .Y(_20995_) );
	NAND2X1 NAND2X1_3636 ( .gnd(gnd), .vdd(vdd), .A(_20995_), .B(_20990_), .Y(_20996_) );
	NOR2X1 NOR2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_20996_), .B(_20986_), .Y(_20997_) );
	AOI22X1 AOI22X1_464 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_11_), .C(registers_r1_11_), .D(_20606__bF_buf3), .Y(_20998_) );
	AOI22X1 AOI22X1_465 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_11_), .C(registers_r5_11_), .D(_20611__bF_buf3), .Y(_20999_) );
	NAND3X1 NAND3X1_3840 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_11_), .B(_20607__bF_buf1), .C(_20574__bF_buf3), .Y(_21000_) );
	OAI21X1 OAI21X1_4709 ( .gnd(gnd), .vdd(vdd), .A(_18045_), .B(_20617__bF_buf3), .C(_21000_), .Y(_21001_) );
	AOI21X1 AOI21X1_3158 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_11_), .B(_20615__bF_buf3), .C(_21001_), .Y(_21002_) );
	NAND3X1 NAND3X1_3841 ( .gnd(gnd), .vdd(vdd), .A(_20998_), .B(_20999_), .C(_21002_), .Y(_21003_) );
	OAI22X1 OAI22X1_500 ( .gnd(gnd), .vdd(vdd), .A(_18051_), .B(_20622__bF_buf3), .C(_18050_), .D(_20621__bF_buf3), .Y(_21004_) );
	OAI22X1 OAI22X1_501 ( .gnd(gnd), .vdd(vdd), .A(_18053_), .B(_20626__bF_buf3), .C(_18054_), .D(_20624__bF_buf3), .Y(_21005_) );
	NOR2X1 NOR2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_21005_), .B(_21004_), .Y(_21006_) );
	OAI22X1 OAI22X1_502 ( .gnd(gnd), .vdd(vdd), .A(_18057_), .B(_20629__bF_buf3), .C(_18058_), .D(_20630__bF_buf3), .Y(_21007_) );
	OAI22X1 OAI22X1_503 ( .gnd(gnd), .vdd(vdd), .A(_18061_), .B(_20633__bF_buf3), .C(_18060_), .D(_20632__bF_buf3), .Y(_21008_) );
	NOR2X1 NOR2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_21007_), .B(_21008_), .Y(_21009_) );
	NAND2X1 NAND2X1_3637 ( .gnd(gnd), .vdd(vdd), .A(_21006_), .B(_21009_), .Y(_21010_) );
	NOR2X1 NOR2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_21003_), .B(_21010_), .Y(_21011_) );
	NAND2X1 NAND2X1_3638 ( .gnd(gnd), .vdd(vdd), .A(_21011_), .B(_20997_), .Y(readB_regOut_11_) );
	NAND3X1 NAND3X1_3842 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_12_), .B(_20559__bF_buf5), .C(_20557__bF_buf6), .Y(_21012_) );
	NAND3X1 NAND3X1_3843 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_12_), .B(_20562__bF_buf5), .C(_20557__bF_buf5), .Y(_21013_) );
	NAND2X1 NAND2X1_3639 ( .gnd(gnd), .vdd(vdd), .A(_21012_), .B(_21013_), .Y(_21014_) );
	OAI22X1 OAI22X1_504 ( .gnd(gnd), .vdd(vdd), .A(_18069_), .B(_20568__bF_buf2), .C(_18070_), .D(_20567__bF_buf2), .Y(_21015_) );
	NOR2X1 NOR2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_21014_), .B(_21015_), .Y(_21016_) );
	OAI22X1 OAI22X1_505 ( .gnd(gnd), .vdd(vdd), .A(_18073_), .B(_20576__bF_buf2), .C(_18074_), .D(_20575__bF_buf2), .Y(_21017_) );
	OAI22X1 OAI22X1_506 ( .gnd(gnd), .vdd(vdd), .A(_18076_), .B(_20581__bF_buf2), .C(_18077_), .D(_20580__bF_buf2), .Y(_21018_) );
	NOR2X1 NOR2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_21018_), .B(_21017_), .Y(_21019_) );
	NAND2X1 NAND2X1_3640 ( .gnd(gnd), .vdd(vdd), .A(_21016_), .B(_21019_), .Y(_21020_) );
	OAI22X1 OAI22X1_507 ( .gnd(gnd), .vdd(vdd), .A(_18082_), .B(_20586__bF_buf2), .C(_18081_), .D(_20585__bF_buf2), .Y(_21021_) );
	NAND3X1 NAND3X1_3844 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_12_), .B(_20588__bF_buf1), .C(_20590__bF_buf7), .Y(_21022_) );
	OAI21X1 OAI21X1_4710 ( .gnd(gnd), .vdd(vdd), .A(_18084_), .B(_20589__bF_buf2), .C(_21022_), .Y(_21023_) );
	NOR2X1 NOR2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_21021_), .B(_21023_), .Y(_21024_) );
	NAND3X1 NAND3X1_3845 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_12_), .B(bLoc_frameOut_4_bF_buf3), .C(_20595__bF_buf2), .Y(_21025_) );
	OAI21X1 OAI21X1_4711 ( .gnd(gnd), .vdd(vdd), .A(_18088_), .B(_20594__bF_buf2), .C(_21025_), .Y(_21026_) );
	NAND3X1 NAND3X1_3846 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_12_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_21027_) );
	OAI21X1 OAI21X1_4712 ( .gnd(gnd), .vdd(vdd), .A(_18091_), .B(_20598__bF_buf2), .C(_21027_), .Y(_21028_) );
	NOR2X1 NOR2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_21026_), .B(_21028_), .Y(_21029_) );
	NAND2X1 NAND2X1_3641 ( .gnd(gnd), .vdd(vdd), .A(_21029_), .B(_21024_), .Y(_21030_) );
	NOR2X1 NOR2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_21030_), .B(_21020_), .Y(_21031_) );
	AOI22X1 AOI22X1_466 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf2), .B(registers_a2_12_), .C(registers_r1_12_), .D(_20606__bF_buf2), .Y(_21032_) );
	AOI22X1 AOI22X1_467 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf2), .B(registers_r4_12_), .C(registers_r5_12_), .D(_20611__bF_buf2), .Y(_21033_) );
	NAND3X1 NAND3X1_3847 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_12_), .B(_20607__bF_buf0), .C(_20574__bF_buf1), .Y(_21034_) );
	OAI21X1 OAI21X1_4713 ( .gnd(gnd), .vdd(vdd), .A(_18099_), .B(_20617__bF_buf2), .C(_21034_), .Y(_21035_) );
	AOI21X1 AOI21X1_3159 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_12_), .B(_20615__bF_buf2), .C(_21035_), .Y(_21036_) );
	NAND3X1 NAND3X1_3848 ( .gnd(gnd), .vdd(vdd), .A(_21032_), .B(_21033_), .C(_21036_), .Y(_21037_) );
	OAI22X1 OAI22X1_508 ( .gnd(gnd), .vdd(vdd), .A(_18105_), .B(_20622__bF_buf2), .C(_18104_), .D(_20621__bF_buf2), .Y(_21038_) );
	OAI22X1 OAI22X1_509 ( .gnd(gnd), .vdd(vdd), .A(_18107_), .B(_20626__bF_buf2), .C(_18108_), .D(_20624__bF_buf2), .Y(_21039_) );
	NOR2X1 NOR2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_21039_), .B(_21038_), .Y(_21040_) );
	OAI22X1 OAI22X1_510 ( .gnd(gnd), .vdd(vdd), .A(_18111_), .B(_20629__bF_buf2), .C(_18112_), .D(_20630__bF_buf2), .Y(_21041_) );
	OAI22X1 OAI22X1_511 ( .gnd(gnd), .vdd(vdd), .A(_18115_), .B(_20633__bF_buf2), .C(_18114_), .D(_20632__bF_buf2), .Y(_21042_) );
	NOR2X1 NOR2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_21041_), .B(_21042_), .Y(_21043_) );
	NAND2X1 NAND2X1_3642 ( .gnd(gnd), .vdd(vdd), .A(_21040_), .B(_21043_), .Y(_21044_) );
	NOR2X1 NOR2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_21037_), .B(_21044_), .Y(_21045_) );
	NAND2X1 NAND2X1_3643 ( .gnd(gnd), .vdd(vdd), .A(_21045_), .B(_21031_), .Y(readB_regOut_12_) );
	NAND3X1 NAND3X1_3849 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_13_), .B(_20559__bF_buf4), .C(_20557__bF_buf4), .Y(_21046_) );
	NAND3X1 NAND3X1_3850 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_13_), .B(_20562__bF_buf4), .C(_20557__bF_buf3), .Y(_21047_) );
	NAND2X1 NAND2X1_3644 ( .gnd(gnd), .vdd(vdd), .A(_21046_), .B(_21047_), .Y(_21048_) );
	OAI22X1 OAI22X1_512 ( .gnd(gnd), .vdd(vdd), .A(_18123_), .B(_20568__bF_buf1), .C(_18124_), .D(_20567__bF_buf1), .Y(_21049_) );
	NOR2X1 NOR2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_21048_), .B(_21049_), .Y(_21050_) );
	OAI22X1 OAI22X1_513 ( .gnd(gnd), .vdd(vdd), .A(_18127_), .B(_20576__bF_buf1), .C(_18128_), .D(_20575__bF_buf1), .Y(_21051_) );
	OAI22X1 OAI22X1_514 ( .gnd(gnd), .vdd(vdd), .A(_18130_), .B(_20581__bF_buf1), .C(_18131_), .D(_20580__bF_buf1), .Y(_21052_) );
	NOR2X1 NOR2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_21052_), .B(_21051_), .Y(_21053_) );
	NAND2X1 NAND2X1_3645 ( .gnd(gnd), .vdd(vdd), .A(_21050_), .B(_21053_), .Y(_21054_) );
	OAI22X1 OAI22X1_515 ( .gnd(gnd), .vdd(vdd), .A(_18136_), .B(_20586__bF_buf1), .C(_18135_), .D(_20585__bF_buf1), .Y(_21055_) );
	NAND3X1 NAND3X1_3851 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_13_), .B(_20588__bF_buf0), .C(_20590__bF_buf5), .Y(_21056_) );
	OAI21X1 OAI21X1_4714 ( .gnd(gnd), .vdd(vdd), .A(_18138_), .B(_20589__bF_buf1), .C(_21056_), .Y(_21057_) );
	NOR2X1 NOR2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_21055_), .B(_21057_), .Y(_21058_) );
	NAND3X1 NAND3X1_3852 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_13_), .B(bLoc_frameOut_4_bF_buf2), .C(_20595__bF_buf1), .Y(_21059_) );
	OAI21X1 OAI21X1_4715 ( .gnd(gnd), .vdd(vdd), .A(_18142_), .B(_20594__bF_buf1), .C(_21059_), .Y(_21060_) );
	NAND3X1 NAND3X1_3853 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_13_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_21061_) );
	OAI21X1 OAI21X1_4716 ( .gnd(gnd), .vdd(vdd), .A(_18145_), .B(_20598__bF_buf1), .C(_21061_), .Y(_21062_) );
	NOR2X1 NOR2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_21060_), .B(_21062_), .Y(_21063_) );
	NAND2X1 NAND2X1_3646 ( .gnd(gnd), .vdd(vdd), .A(_21063_), .B(_21058_), .Y(_21064_) );
	NOR2X1 NOR2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_21064_), .B(_21054_), .Y(_21065_) );
	AOI22X1 AOI22X1_468 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf1), .B(registers_a2_13_), .C(registers_r1_13_), .D(_20606__bF_buf1), .Y(_21066_) );
	AOI22X1 AOI22X1_469 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf1), .B(registers_r4_13_), .C(registers_r5_13_), .D(_20611__bF_buf1), .Y(_21067_) );
	NAND3X1 NAND3X1_3854 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_13_), .B(_20607__bF_buf4), .C(_20574__bF_buf7), .Y(_21068_) );
	OAI21X1 OAI21X1_4717 ( .gnd(gnd), .vdd(vdd), .A(_18153_), .B(_20617__bF_buf1), .C(_21068_), .Y(_21069_) );
	AOI21X1 AOI21X1_3160 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_13_), .B(_20615__bF_buf1), .C(_21069_), .Y(_21070_) );
	NAND3X1 NAND3X1_3855 ( .gnd(gnd), .vdd(vdd), .A(_21066_), .B(_21067_), .C(_21070_), .Y(_21071_) );
	OAI22X1 OAI22X1_516 ( .gnd(gnd), .vdd(vdd), .A(_18159_), .B(_20622__bF_buf1), .C(_18158_), .D(_20621__bF_buf1), .Y(_21072_) );
	OAI22X1 OAI22X1_517 ( .gnd(gnd), .vdd(vdd), .A(_18161_), .B(_20626__bF_buf1), .C(_18162_), .D(_20624__bF_buf1), .Y(_21073_) );
	NOR2X1 NOR2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_21073_), .B(_21072_), .Y(_21074_) );
	OAI22X1 OAI22X1_518 ( .gnd(gnd), .vdd(vdd), .A(_18165_), .B(_20629__bF_buf1), .C(_18166_), .D(_20630__bF_buf1), .Y(_21075_) );
	OAI22X1 OAI22X1_519 ( .gnd(gnd), .vdd(vdd), .A(_18169_), .B(_20633__bF_buf1), .C(_18168_), .D(_20632__bF_buf1), .Y(_21076_) );
	NOR2X1 NOR2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_21075_), .B(_21076_), .Y(_21077_) );
	NAND2X1 NAND2X1_3647 ( .gnd(gnd), .vdd(vdd), .A(_21074_), .B(_21077_), .Y(_21078_) );
	NOR2X1 NOR2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_21071_), .B(_21078_), .Y(_21079_) );
	NAND2X1 NAND2X1_3648 ( .gnd(gnd), .vdd(vdd), .A(_21079_), .B(_21065_), .Y(readB_regOut_13_) );
	NAND3X1 NAND3X1_3856 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_14_), .B(_20559__bF_buf3), .C(_20557__bF_buf2), .Y(_21080_) );
	NAND3X1 NAND3X1_3857 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_14_), .B(_20562__bF_buf3), .C(_20557__bF_buf1), .Y(_21081_) );
	NAND2X1 NAND2X1_3649 ( .gnd(gnd), .vdd(vdd), .A(_21080_), .B(_21081_), .Y(_21082_) );
	OAI22X1 OAI22X1_520 ( .gnd(gnd), .vdd(vdd), .A(_18177_), .B(_20568__bF_buf0), .C(_18178_), .D(_20567__bF_buf0), .Y(_21083_) );
	NOR2X1 NOR2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_21082_), .B(_21083_), .Y(_21084_) );
	OAI22X1 OAI22X1_521 ( .gnd(gnd), .vdd(vdd), .A(_18181_), .B(_20576__bF_buf0), .C(_18182_), .D(_20575__bF_buf0), .Y(_21085_) );
	OAI22X1 OAI22X1_522 ( .gnd(gnd), .vdd(vdd), .A(_18184_), .B(_20581__bF_buf0), .C(_18185_), .D(_20580__bF_buf0), .Y(_21086_) );
	NOR2X1 NOR2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_21086_), .B(_21085_), .Y(_21087_) );
	NAND2X1 NAND2X1_3650 ( .gnd(gnd), .vdd(vdd), .A(_21084_), .B(_21087_), .Y(_21088_) );
	OAI22X1 OAI22X1_523 ( .gnd(gnd), .vdd(vdd), .A(_18190_), .B(_20586__bF_buf0), .C(_18189_), .D(_20585__bF_buf0), .Y(_21089_) );
	NAND3X1 NAND3X1_3858 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_14_), .B(_20588__bF_buf5), .C(_20590__bF_buf3), .Y(_21090_) );
	OAI21X1 OAI21X1_4718 ( .gnd(gnd), .vdd(vdd), .A(_18192_), .B(_20589__bF_buf0), .C(_21090_), .Y(_21091_) );
	NOR2X1 NOR2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_21089_), .B(_21091_), .Y(_21092_) );
	NAND3X1 NAND3X1_3859 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_14_), .B(bLoc_frameOut_4_bF_buf1), .C(_20595__bF_buf0), .Y(_21093_) );
	OAI21X1 OAI21X1_4719 ( .gnd(gnd), .vdd(vdd), .A(_18196_), .B(_20594__bF_buf0), .C(_21093_), .Y(_21094_) );
	NAND3X1 NAND3X1_3860 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_14_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_21095_) );
	OAI21X1 OAI21X1_4720 ( .gnd(gnd), .vdd(vdd), .A(_18199_), .B(_20598__bF_buf0), .C(_21095_), .Y(_21096_) );
	NOR2X1 NOR2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_21094_), .B(_21096_), .Y(_21097_) );
	NAND2X1 NAND2X1_3651 ( .gnd(gnd), .vdd(vdd), .A(_21097_), .B(_21092_), .Y(_21098_) );
	NOR2X1 NOR2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_21098_), .B(_21088_), .Y(_21099_) );
	AOI22X1 AOI22X1_470 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf0), .B(registers_a2_14_), .C(registers_r1_14_), .D(_20606__bF_buf0), .Y(_21100_) );
	AOI22X1 AOI22X1_471 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf0), .B(registers_r4_14_), .C(registers_r5_14_), .D(_20611__bF_buf0), .Y(_21101_) );
	NAND3X1 NAND3X1_3861 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_14_), .B(_20607__bF_buf3), .C(_20574__bF_buf5), .Y(_21102_) );
	OAI21X1 OAI21X1_4721 ( .gnd(gnd), .vdd(vdd), .A(_18207_), .B(_20617__bF_buf0), .C(_21102_), .Y(_21103_) );
	AOI21X1 AOI21X1_3161 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_14_), .B(_20615__bF_buf0), .C(_21103_), .Y(_21104_) );
	NAND3X1 NAND3X1_3862 ( .gnd(gnd), .vdd(vdd), .A(_21100_), .B(_21101_), .C(_21104_), .Y(_21105_) );
	OAI22X1 OAI22X1_524 ( .gnd(gnd), .vdd(vdd), .A(_18213_), .B(_20622__bF_buf0), .C(_18212_), .D(_20621__bF_buf0), .Y(_21106_) );
	OAI22X1 OAI22X1_525 ( .gnd(gnd), .vdd(vdd), .A(_18215_), .B(_20626__bF_buf0), .C(_18216_), .D(_20624__bF_buf0), .Y(_21107_) );
	NOR2X1 NOR2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_21107_), .B(_21106_), .Y(_21108_) );
	OAI22X1 OAI22X1_526 ( .gnd(gnd), .vdd(vdd), .A(_18219_), .B(_20629__bF_buf0), .C(_18220_), .D(_20630__bF_buf0), .Y(_21109_) );
	OAI22X1 OAI22X1_527 ( .gnd(gnd), .vdd(vdd), .A(_18223_), .B(_20633__bF_buf0), .C(_18222_), .D(_20632__bF_buf0), .Y(_21110_) );
	NOR2X1 NOR2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_21109_), .B(_21110_), .Y(_21111_) );
	NAND2X1 NAND2X1_3652 ( .gnd(gnd), .vdd(vdd), .A(_21108_), .B(_21111_), .Y(_21112_) );
	NOR2X1 NOR2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_21105_), .B(_21112_), .Y(_21113_) );
	NAND2X1 NAND2X1_3653 ( .gnd(gnd), .vdd(vdd), .A(_21113_), .B(_21099_), .Y(readB_regOut_14_) );
	NAND3X1 NAND3X1_3863 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_15_), .B(_20559__bF_buf2), .C(_20557__bF_buf0), .Y(_21114_) );
	NAND3X1 NAND3X1_3864 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_15_), .B(_20562__bF_buf2), .C(_20557__bF_buf7), .Y(_21115_) );
	NAND2X1 NAND2X1_3654 ( .gnd(gnd), .vdd(vdd), .A(_21114_), .B(_21115_), .Y(_21116_) );
	OAI22X1 OAI22X1_528 ( .gnd(gnd), .vdd(vdd), .A(_18231_), .B(_20568__bF_buf4), .C(_18232_), .D(_20567__bF_buf4), .Y(_21117_) );
	NOR2X1 NOR2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_21116_), .B(_21117_), .Y(_21118_) );
	OAI22X1 OAI22X1_529 ( .gnd(gnd), .vdd(vdd), .A(_18235_), .B(_20576__bF_buf4), .C(_18236_), .D(_20575__bF_buf4), .Y(_21119_) );
	OAI22X1 OAI22X1_530 ( .gnd(gnd), .vdd(vdd), .A(_18238_), .B(_20581__bF_buf4), .C(_18239_), .D(_20580__bF_buf4), .Y(_21120_) );
	NOR2X1 NOR2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_21120_), .B(_21119_), .Y(_21121_) );
	NAND2X1 NAND2X1_3655 ( .gnd(gnd), .vdd(vdd), .A(_21118_), .B(_21121_), .Y(_21122_) );
	OAI22X1 OAI22X1_531 ( .gnd(gnd), .vdd(vdd), .A(_18244_), .B(_20586__bF_buf4), .C(_18243_), .D(_20585__bF_buf4), .Y(_21123_) );
	NAND3X1 NAND3X1_3865 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_15_), .B(_20588__bF_buf4), .C(_20590__bF_buf1), .Y(_21124_) );
	OAI21X1 OAI21X1_4722 ( .gnd(gnd), .vdd(vdd), .A(_18246_), .B(_20589__bF_buf4), .C(_21124_), .Y(_21125_) );
	NOR2X1 NOR2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_21123_), .B(_21125_), .Y(_21126_) );
	NAND3X1 NAND3X1_3866 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_15_), .B(bLoc_frameOut_4_bF_buf0), .C(_20595__bF_buf4), .Y(_21127_) );
	OAI21X1 OAI21X1_4723 ( .gnd(gnd), .vdd(vdd), .A(_18250_), .B(_20594__bF_buf4), .C(_21127_), .Y(_21128_) );
	NAND3X1 NAND3X1_3867 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_15_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_21129_) );
	OAI21X1 OAI21X1_4724 ( .gnd(gnd), .vdd(vdd), .A(_18253_), .B(_20598__bF_buf4), .C(_21129_), .Y(_21130_) );
	NOR2X1 NOR2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_21128_), .B(_21130_), .Y(_21131_) );
	NAND2X1 NAND2X1_3656 ( .gnd(gnd), .vdd(vdd), .A(_21131_), .B(_21126_), .Y(_21132_) );
	NOR2X1 NOR2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_21132_), .B(_21122_), .Y(_21133_) );
	AOI22X1 AOI22X1_472 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_15_), .C(registers_r1_15_), .D(_20606__bF_buf4), .Y(_21134_) );
	AOI22X1 AOI22X1_473 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_15_), .C(registers_r5_15_), .D(_20611__bF_buf4), .Y(_21135_) );
	NAND3X1 NAND3X1_3868 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_15_), .B(_20607__bF_buf2), .C(_20574__bF_buf3), .Y(_21136_) );
	OAI21X1 OAI21X1_4725 ( .gnd(gnd), .vdd(vdd), .A(_18261_), .B(_20617__bF_buf4), .C(_21136_), .Y(_21137_) );
	AOI21X1 AOI21X1_3162 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_15_), .B(_20615__bF_buf4), .C(_21137_), .Y(_21138_) );
	NAND3X1 NAND3X1_3869 ( .gnd(gnd), .vdd(vdd), .A(_21134_), .B(_21135_), .C(_21138_), .Y(_21139_) );
	OAI22X1 OAI22X1_532 ( .gnd(gnd), .vdd(vdd), .A(_18267_), .B(_20622__bF_buf4), .C(_18266_), .D(_20621__bF_buf4), .Y(_21140_) );
	OAI22X1 OAI22X1_533 ( .gnd(gnd), .vdd(vdd), .A(_18269_), .B(_20626__bF_buf4), .C(_18270_), .D(_20624__bF_buf4), .Y(_21141_) );
	NOR2X1 NOR2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_21141_), .B(_21140_), .Y(_21142_) );
	OAI22X1 OAI22X1_534 ( .gnd(gnd), .vdd(vdd), .A(_18273_), .B(_20629__bF_buf4), .C(_18274_), .D(_20630__bF_buf4), .Y(_21143_) );
	OAI22X1 OAI22X1_535 ( .gnd(gnd), .vdd(vdd), .A(_18277_), .B(_20633__bF_buf4), .C(_18276_), .D(_20632__bF_buf4), .Y(_21144_) );
	NOR2X1 NOR2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_21143_), .B(_21144_), .Y(_21145_) );
	NAND2X1 NAND2X1_3657 ( .gnd(gnd), .vdd(vdd), .A(_21142_), .B(_21145_), .Y(_21146_) );
	NOR2X1 NOR2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_21139_), .B(_21146_), .Y(_21147_) );
	NAND2X1 NAND2X1_3658 ( .gnd(gnd), .vdd(vdd), .A(_21147_), .B(_21133_), .Y(readB_regOut_15_) );
	NAND3X1 NAND3X1_3870 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_16_), .B(_20559__bF_buf1), .C(_20557__bF_buf6), .Y(_21148_) );
	NAND3X1 NAND3X1_3871 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_16_), .B(_20562__bF_buf1), .C(_20557__bF_buf5), .Y(_21149_) );
	NAND2X1 NAND2X1_3659 ( .gnd(gnd), .vdd(vdd), .A(_21148_), .B(_21149_), .Y(_21150_) );
	OAI22X1 OAI22X1_536 ( .gnd(gnd), .vdd(vdd), .A(_18285_), .B(_20568__bF_buf3), .C(_18286_), .D(_20567__bF_buf3), .Y(_21151_) );
	NOR2X1 NOR2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_21150_), .B(_21151_), .Y(_21152_) );
	OAI22X1 OAI22X1_537 ( .gnd(gnd), .vdd(vdd), .A(_18289_), .B(_20576__bF_buf3), .C(_18290_), .D(_20575__bF_buf3), .Y(_21153_) );
	OAI22X1 OAI22X1_538 ( .gnd(gnd), .vdd(vdd), .A(_18292_), .B(_20581__bF_buf3), .C(_18293_), .D(_20580__bF_buf3), .Y(_21154_) );
	NOR2X1 NOR2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_21154_), .B(_21153_), .Y(_21155_) );
	NAND2X1 NAND2X1_3660 ( .gnd(gnd), .vdd(vdd), .A(_21152_), .B(_21155_), .Y(_21156_) );
	OAI22X1 OAI22X1_539 ( .gnd(gnd), .vdd(vdd), .A(_18298_), .B(_20586__bF_buf3), .C(_18297_), .D(_20585__bF_buf3), .Y(_21157_) );
	NAND3X1 NAND3X1_3872 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_16_), .B(_20588__bF_buf3), .C(_20590__bF_buf7), .Y(_21158_) );
	OAI21X1 OAI21X1_4726 ( .gnd(gnd), .vdd(vdd), .A(_18300_), .B(_20589__bF_buf3), .C(_21158_), .Y(_21159_) );
	NOR2X1 NOR2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_21157_), .B(_21159_), .Y(_21160_) );
	NAND3X1 NAND3X1_3873 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_16_), .B(bLoc_frameOut_4_bF_buf6), .C(_20595__bF_buf3), .Y(_21161_) );
	OAI21X1 OAI21X1_4727 ( .gnd(gnd), .vdd(vdd), .A(_18304_), .B(_20594__bF_buf3), .C(_21161_), .Y(_21162_) );
	NAND3X1 NAND3X1_3874 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_16_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_21163_) );
	OAI21X1 OAI21X1_4728 ( .gnd(gnd), .vdd(vdd), .A(_18307_), .B(_20598__bF_buf3), .C(_21163_), .Y(_21164_) );
	NOR2X1 NOR2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_21162_), .B(_21164_), .Y(_21165_) );
	NAND2X1 NAND2X1_3661 ( .gnd(gnd), .vdd(vdd), .A(_21165_), .B(_21160_), .Y(_21166_) );
	NOR2X1 NOR2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_21166_), .B(_21156_), .Y(_21167_) );
	AOI22X1 AOI22X1_474 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_16_), .C(registers_r1_16_), .D(_20606__bF_buf3), .Y(_21168_) );
	AOI22X1 AOI22X1_475 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_16_), .C(registers_r5_16_), .D(_20611__bF_buf3), .Y(_21169_) );
	NAND3X1 NAND3X1_3875 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_16_), .B(_20607__bF_buf1), .C(_20574__bF_buf1), .Y(_21170_) );
	OAI21X1 OAI21X1_4729 ( .gnd(gnd), .vdd(vdd), .A(_18315_), .B(_20617__bF_buf3), .C(_21170_), .Y(_21171_) );
	AOI21X1 AOI21X1_3163 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_16_), .B(_20615__bF_buf3), .C(_21171_), .Y(_21172_) );
	NAND3X1 NAND3X1_3876 ( .gnd(gnd), .vdd(vdd), .A(_21168_), .B(_21169_), .C(_21172_), .Y(_21173_) );
	OAI22X1 OAI22X1_540 ( .gnd(gnd), .vdd(vdd), .A(_18321_), .B(_20622__bF_buf3), .C(_18320_), .D(_20621__bF_buf3), .Y(_21174_) );
	OAI22X1 OAI22X1_541 ( .gnd(gnd), .vdd(vdd), .A(_18323_), .B(_20626__bF_buf3), .C(_18324_), .D(_20624__bF_buf3), .Y(_21175_) );
	NOR2X1 NOR2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_21175_), .B(_21174_), .Y(_21176_) );
	OAI22X1 OAI22X1_542 ( .gnd(gnd), .vdd(vdd), .A(_18327_), .B(_20629__bF_buf3), .C(_18328_), .D(_20630__bF_buf3), .Y(_21177_) );
	OAI22X1 OAI22X1_543 ( .gnd(gnd), .vdd(vdd), .A(_18331_), .B(_20633__bF_buf3), .C(_18330_), .D(_20632__bF_buf3), .Y(_21178_) );
	NOR2X1 NOR2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_21177_), .B(_21178_), .Y(_21179_) );
	NAND2X1 NAND2X1_3662 ( .gnd(gnd), .vdd(vdd), .A(_21176_), .B(_21179_), .Y(_21180_) );
	NOR2X1 NOR2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_21173_), .B(_21180_), .Y(_21181_) );
	NAND2X1 NAND2X1_3663 ( .gnd(gnd), .vdd(vdd), .A(_21181_), .B(_21167_), .Y(readB_regOut_16_) );
	NAND3X1 NAND3X1_3877 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_17_), .B(_20559__bF_buf0), .C(_20557__bF_buf4), .Y(_21182_) );
	NAND3X1 NAND3X1_3878 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_17_), .B(_20562__bF_buf0), .C(_20557__bF_buf3), .Y(_21183_) );
	NAND2X1 NAND2X1_3664 ( .gnd(gnd), .vdd(vdd), .A(_21182_), .B(_21183_), .Y(_21184_) );
	OAI22X1 OAI22X1_544 ( .gnd(gnd), .vdd(vdd), .A(_18339_), .B(_20568__bF_buf2), .C(_18340_), .D(_20567__bF_buf2), .Y(_21185_) );
	NOR2X1 NOR2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_21184_), .B(_21185_), .Y(_21186_) );
	OAI22X1 OAI22X1_545 ( .gnd(gnd), .vdd(vdd), .A(_18343_), .B(_20576__bF_buf2), .C(_18344_), .D(_20575__bF_buf2), .Y(_21187_) );
	OAI22X1 OAI22X1_546 ( .gnd(gnd), .vdd(vdd), .A(_18346_), .B(_20581__bF_buf2), .C(_18347_), .D(_20580__bF_buf2), .Y(_21188_) );
	NOR2X1 NOR2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_21188_), .B(_21187_), .Y(_21189_) );
	NAND2X1 NAND2X1_3665 ( .gnd(gnd), .vdd(vdd), .A(_21186_), .B(_21189_), .Y(_21190_) );
	OAI22X1 OAI22X1_547 ( .gnd(gnd), .vdd(vdd), .A(_18352_), .B(_20586__bF_buf2), .C(_18351_), .D(_20585__bF_buf2), .Y(_21191_) );
	NAND3X1 NAND3X1_3879 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_17_), .B(_20588__bF_buf2), .C(_20590__bF_buf5), .Y(_21192_) );
	OAI21X1 OAI21X1_4730 ( .gnd(gnd), .vdd(vdd), .A(_18354_), .B(_20589__bF_buf2), .C(_21192_), .Y(_21193_) );
	NOR2X1 NOR2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_21191_), .B(_21193_), .Y(_21194_) );
	NAND3X1 NAND3X1_3880 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_17_), .B(bLoc_frameOut_4_bF_buf5), .C(_20595__bF_buf2), .Y(_21195_) );
	OAI21X1 OAI21X1_4731 ( .gnd(gnd), .vdd(vdd), .A(_18358_), .B(_20594__bF_buf2), .C(_21195_), .Y(_21196_) );
	NAND3X1 NAND3X1_3881 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_17_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_21197_) );
	OAI21X1 OAI21X1_4732 ( .gnd(gnd), .vdd(vdd), .A(_18361_), .B(_20598__bF_buf2), .C(_21197_), .Y(_21198_) );
	NOR2X1 NOR2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_21196_), .B(_21198_), .Y(_21199_) );
	NAND2X1 NAND2X1_3666 ( .gnd(gnd), .vdd(vdd), .A(_21199_), .B(_21194_), .Y(_21200_) );
	NOR2X1 NOR2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_21200_), .B(_21190_), .Y(_21201_) );
	AOI22X1 AOI22X1_476 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf2), .B(registers_a2_17_), .C(registers_r1_17_), .D(_20606__bF_buf2), .Y(_21202_) );
	AOI22X1 AOI22X1_477 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf2), .B(registers_r4_17_), .C(registers_r5_17_), .D(_20611__bF_buf2), .Y(_21203_) );
	NAND3X1 NAND3X1_3882 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_17_), .B(_20607__bF_buf0), .C(_20574__bF_buf7), .Y(_21204_) );
	OAI21X1 OAI21X1_4733 ( .gnd(gnd), .vdd(vdd), .A(_18369_), .B(_20617__bF_buf2), .C(_21204_), .Y(_21205_) );
	AOI21X1 AOI21X1_3164 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_17_), .B(_20615__bF_buf2), .C(_21205_), .Y(_21206_) );
	NAND3X1 NAND3X1_3883 ( .gnd(gnd), .vdd(vdd), .A(_21202_), .B(_21203_), .C(_21206_), .Y(_21207_) );
	OAI22X1 OAI22X1_548 ( .gnd(gnd), .vdd(vdd), .A(_18375_), .B(_20622__bF_buf2), .C(_18374_), .D(_20621__bF_buf2), .Y(_21208_) );
	OAI22X1 OAI22X1_549 ( .gnd(gnd), .vdd(vdd), .A(_18377_), .B(_20626__bF_buf2), .C(_18378_), .D(_20624__bF_buf2), .Y(_21209_) );
	NOR2X1 NOR2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_21209_), .B(_21208_), .Y(_21210_) );
	OAI22X1 OAI22X1_550 ( .gnd(gnd), .vdd(vdd), .A(_18381_), .B(_20629__bF_buf2), .C(_18382_), .D(_20630__bF_buf2), .Y(_21211_) );
	OAI22X1 OAI22X1_551 ( .gnd(gnd), .vdd(vdd), .A(_18385_), .B(_20633__bF_buf2), .C(_18384_), .D(_20632__bF_buf2), .Y(_21212_) );
	NOR2X1 NOR2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_21211_), .B(_21212_), .Y(_21213_) );
	NAND2X1 NAND2X1_3667 ( .gnd(gnd), .vdd(vdd), .A(_21210_), .B(_21213_), .Y(_21214_) );
	NOR2X1 NOR2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_21207_), .B(_21214_), .Y(_21215_) );
	NAND2X1 NAND2X1_3668 ( .gnd(gnd), .vdd(vdd), .A(_21215_), .B(_21201_), .Y(readB_regOut_17_) );
	NAND3X1 NAND3X1_3884 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_18_), .B(_20559__bF_buf5), .C(_20557__bF_buf2), .Y(_21216_) );
	NAND3X1 NAND3X1_3885 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_18_), .B(_20562__bF_buf5), .C(_20557__bF_buf1), .Y(_21217_) );
	NAND2X1 NAND2X1_3669 ( .gnd(gnd), .vdd(vdd), .A(_21216_), .B(_21217_), .Y(_21218_) );
	OAI22X1 OAI22X1_552 ( .gnd(gnd), .vdd(vdd), .A(_18393_), .B(_20568__bF_buf1), .C(_18394_), .D(_20567__bF_buf1), .Y(_21219_) );
	NOR2X1 NOR2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_21218_), .B(_21219_), .Y(_21220_) );
	OAI22X1 OAI22X1_553 ( .gnd(gnd), .vdd(vdd), .A(_18397_), .B(_20576__bF_buf1), .C(_18398_), .D(_20575__bF_buf1), .Y(_21221_) );
	OAI22X1 OAI22X1_554 ( .gnd(gnd), .vdd(vdd), .A(_18400_), .B(_20581__bF_buf1), .C(_18401_), .D(_20580__bF_buf1), .Y(_21222_) );
	NOR2X1 NOR2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_21222_), .B(_21221_), .Y(_21223_) );
	NAND2X1 NAND2X1_3670 ( .gnd(gnd), .vdd(vdd), .A(_21220_), .B(_21223_), .Y(_21224_) );
	OAI22X1 OAI22X1_555 ( .gnd(gnd), .vdd(vdd), .A(_18406_), .B(_20586__bF_buf1), .C(_18405_), .D(_20585__bF_buf1), .Y(_21225_) );
	NAND3X1 NAND3X1_3886 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_18_), .B(_20588__bF_buf1), .C(_20590__bF_buf3), .Y(_21226_) );
	OAI21X1 OAI21X1_4734 ( .gnd(gnd), .vdd(vdd), .A(_18408_), .B(_20589__bF_buf1), .C(_21226_), .Y(_21227_) );
	NOR2X1 NOR2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_21225_), .B(_21227_), .Y(_21228_) );
	NAND3X1 NAND3X1_3887 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_18_), .B(bLoc_frameOut_4_bF_buf4), .C(_20595__bF_buf1), .Y(_21229_) );
	OAI21X1 OAI21X1_4735 ( .gnd(gnd), .vdd(vdd), .A(_18412_), .B(_20594__bF_buf1), .C(_21229_), .Y(_21230_) );
	NAND3X1 NAND3X1_3888 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_18_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_21231_) );
	OAI21X1 OAI21X1_4736 ( .gnd(gnd), .vdd(vdd), .A(_18415_), .B(_20598__bF_buf1), .C(_21231_), .Y(_21232_) );
	NOR2X1 NOR2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_21230_), .B(_21232_), .Y(_21233_) );
	NAND2X1 NAND2X1_3671 ( .gnd(gnd), .vdd(vdd), .A(_21233_), .B(_21228_), .Y(_21234_) );
	NOR2X1 NOR2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_21234_), .B(_21224_), .Y(_21235_) );
	AOI22X1 AOI22X1_478 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf1), .B(registers_a2_18_), .C(registers_r1_18_), .D(_20606__bF_buf1), .Y(_21236_) );
	AOI22X1 AOI22X1_479 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf1), .B(registers_r4_18_), .C(registers_r5_18_), .D(_20611__bF_buf1), .Y(_21237_) );
	NAND3X1 NAND3X1_3889 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_18_), .B(_20607__bF_buf4), .C(_20574__bF_buf5), .Y(_21238_) );
	OAI21X1 OAI21X1_4737 ( .gnd(gnd), .vdd(vdd), .A(_18423_), .B(_20617__bF_buf1), .C(_21238_), .Y(_21239_) );
	AOI21X1 AOI21X1_3165 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_18_), .B(_20615__bF_buf1), .C(_21239_), .Y(_21240_) );
	NAND3X1 NAND3X1_3890 ( .gnd(gnd), .vdd(vdd), .A(_21236_), .B(_21237_), .C(_21240_), .Y(_21241_) );
	OAI22X1 OAI22X1_556 ( .gnd(gnd), .vdd(vdd), .A(_18429_), .B(_20622__bF_buf1), .C(_18428_), .D(_20621__bF_buf1), .Y(_21242_) );
	OAI22X1 OAI22X1_557 ( .gnd(gnd), .vdd(vdd), .A(_18431_), .B(_20626__bF_buf1), .C(_18432_), .D(_20624__bF_buf1), .Y(_21243_) );
	NOR2X1 NOR2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_21243_), .B(_21242_), .Y(_21244_) );
	OAI22X1 OAI22X1_558 ( .gnd(gnd), .vdd(vdd), .A(_18435_), .B(_20629__bF_buf1), .C(_18436_), .D(_20630__bF_buf1), .Y(_21245_) );
	OAI22X1 OAI22X1_559 ( .gnd(gnd), .vdd(vdd), .A(_18439_), .B(_20633__bF_buf1), .C(_18438_), .D(_20632__bF_buf1), .Y(_21246_) );
	NOR2X1 NOR2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_21245_), .B(_21246_), .Y(_21247_) );
	NAND2X1 NAND2X1_3672 ( .gnd(gnd), .vdd(vdd), .A(_21244_), .B(_21247_), .Y(_21248_) );
	NOR2X1 NOR2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_21241_), .B(_21248_), .Y(_21249_) );
	NAND2X1 NAND2X1_3673 ( .gnd(gnd), .vdd(vdd), .A(_21249_), .B(_21235_), .Y(readB_regOut_18_) );
	NAND3X1 NAND3X1_3891 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_19_), .B(_20559__bF_buf4), .C(_20557__bF_buf0), .Y(_21250_) );
	NAND3X1 NAND3X1_3892 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_19_), .B(_20562__bF_buf4), .C(_20557__bF_buf7), .Y(_21251_) );
	NAND2X1 NAND2X1_3674 ( .gnd(gnd), .vdd(vdd), .A(_21250_), .B(_21251_), .Y(_21252_) );
	OAI22X1 OAI22X1_560 ( .gnd(gnd), .vdd(vdd), .A(_18447_), .B(_20568__bF_buf0), .C(_18448_), .D(_20567__bF_buf0), .Y(_21253_) );
	NOR2X1 NOR2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_21252_), .B(_21253_), .Y(_21254_) );
	OAI22X1 OAI22X1_561 ( .gnd(gnd), .vdd(vdd), .A(_18451_), .B(_20576__bF_buf0), .C(_18452_), .D(_20575__bF_buf0), .Y(_21255_) );
	OAI22X1 OAI22X1_562 ( .gnd(gnd), .vdd(vdd), .A(_18454_), .B(_20581__bF_buf0), .C(_18455_), .D(_20580__bF_buf0), .Y(_21256_) );
	NOR2X1 NOR2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_21256_), .B(_21255_), .Y(_21257_) );
	NAND2X1 NAND2X1_3675 ( .gnd(gnd), .vdd(vdd), .A(_21254_), .B(_21257_), .Y(_21258_) );
	OAI22X1 OAI22X1_563 ( .gnd(gnd), .vdd(vdd), .A(_18460_), .B(_20586__bF_buf0), .C(_18459_), .D(_20585__bF_buf0), .Y(_21259_) );
	NAND3X1 NAND3X1_3893 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_19_), .B(_20588__bF_buf0), .C(_20590__bF_buf1), .Y(_21260_) );
	OAI21X1 OAI21X1_4738 ( .gnd(gnd), .vdd(vdd), .A(_18462_), .B(_20589__bF_buf0), .C(_21260_), .Y(_21261_) );
	NOR2X1 NOR2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_21259_), .B(_21261_), .Y(_21262_) );
	NAND3X1 NAND3X1_3894 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_19_), .B(bLoc_frameOut_4_bF_buf3), .C(_20595__bF_buf0), .Y(_21263_) );
	OAI21X1 OAI21X1_4739 ( .gnd(gnd), .vdd(vdd), .A(_18466_), .B(_20594__bF_buf0), .C(_21263_), .Y(_21264_) );
	NAND3X1 NAND3X1_3895 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_19_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_21265_) );
	OAI21X1 OAI21X1_4740 ( .gnd(gnd), .vdd(vdd), .A(_18469_), .B(_20598__bF_buf0), .C(_21265_), .Y(_21266_) );
	NOR2X1 NOR2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_21264_), .B(_21266_), .Y(_21267_) );
	NAND2X1 NAND2X1_3676 ( .gnd(gnd), .vdd(vdd), .A(_21267_), .B(_21262_), .Y(_21268_) );
	NOR2X1 NOR2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_21268_), .B(_21258_), .Y(_21269_) );
	AOI22X1 AOI22X1_480 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf0), .B(registers_a2_19_), .C(registers_r1_19_), .D(_20606__bF_buf0), .Y(_21270_) );
	AOI22X1 AOI22X1_481 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf0), .B(registers_r4_19_), .C(registers_r5_19_), .D(_20611__bF_buf0), .Y(_21271_) );
	NAND3X1 NAND3X1_3896 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_19_), .B(_20607__bF_buf3), .C(_20574__bF_buf3), .Y(_21272_) );
	OAI21X1 OAI21X1_4741 ( .gnd(gnd), .vdd(vdd), .A(_18477_), .B(_20617__bF_buf0), .C(_21272_), .Y(_21273_) );
	AOI21X1 AOI21X1_3166 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_19_), .B(_20615__bF_buf0), .C(_21273_), .Y(_21274_) );
	NAND3X1 NAND3X1_3897 ( .gnd(gnd), .vdd(vdd), .A(_21270_), .B(_21271_), .C(_21274_), .Y(_21275_) );
	OAI22X1 OAI22X1_564 ( .gnd(gnd), .vdd(vdd), .A(_18483_), .B(_20622__bF_buf0), .C(_18482_), .D(_20621__bF_buf0), .Y(_21276_) );
	OAI22X1 OAI22X1_565 ( .gnd(gnd), .vdd(vdd), .A(_18485_), .B(_20626__bF_buf0), .C(_18486_), .D(_20624__bF_buf0), .Y(_21277_) );
	NOR2X1 NOR2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_21277_), .B(_21276_), .Y(_21278_) );
	OAI22X1 OAI22X1_566 ( .gnd(gnd), .vdd(vdd), .A(_18489_), .B(_20629__bF_buf0), .C(_18490_), .D(_20630__bF_buf0), .Y(_21279_) );
	OAI22X1 OAI22X1_567 ( .gnd(gnd), .vdd(vdd), .A(_18493_), .B(_20633__bF_buf0), .C(_18492_), .D(_20632__bF_buf0), .Y(_21280_) );
	NOR2X1 NOR2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_21279_), .B(_21280_), .Y(_21281_) );
	NAND2X1 NAND2X1_3677 ( .gnd(gnd), .vdd(vdd), .A(_21278_), .B(_21281_), .Y(_21282_) );
	NOR2X1 NOR2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_21275_), .B(_21282_), .Y(_21283_) );
	NAND2X1 NAND2X1_3678 ( .gnd(gnd), .vdd(vdd), .A(_21283_), .B(_21269_), .Y(readB_regOut_19_) );
	NAND3X1 NAND3X1_3898 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_20_), .B(_20559__bF_buf3), .C(_20557__bF_buf6), .Y(_21284_) );
	NAND3X1 NAND3X1_3899 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_20_), .B(_20562__bF_buf3), .C(_20557__bF_buf5), .Y(_21285_) );
	NAND2X1 NAND2X1_3679 ( .gnd(gnd), .vdd(vdd), .A(_21284_), .B(_21285_), .Y(_21286_) );
	OAI22X1 OAI22X1_568 ( .gnd(gnd), .vdd(vdd), .A(_18501_), .B(_20568__bF_buf4), .C(_18502_), .D(_20567__bF_buf4), .Y(_21287_) );
	NOR2X1 NOR2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_21286_), .B(_21287_), .Y(_21288_) );
	OAI22X1 OAI22X1_569 ( .gnd(gnd), .vdd(vdd), .A(_18505_), .B(_20576__bF_buf4), .C(_18506_), .D(_20575__bF_buf4), .Y(_21289_) );
	OAI22X1 OAI22X1_570 ( .gnd(gnd), .vdd(vdd), .A(_18508_), .B(_20581__bF_buf4), .C(_18509_), .D(_20580__bF_buf4), .Y(_21290_) );
	NOR2X1 NOR2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_21290_), .B(_21289_), .Y(_21291_) );
	NAND2X1 NAND2X1_3680 ( .gnd(gnd), .vdd(vdd), .A(_21288_), .B(_21291_), .Y(_21292_) );
	OAI22X1 OAI22X1_571 ( .gnd(gnd), .vdd(vdd), .A(_18514_), .B(_20586__bF_buf4), .C(_18513_), .D(_20585__bF_buf4), .Y(_21293_) );
	NAND3X1 NAND3X1_3900 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_20_), .B(_20588__bF_buf5), .C(_20590__bF_buf7), .Y(_21294_) );
	OAI21X1 OAI21X1_4742 ( .gnd(gnd), .vdd(vdd), .A(_18516_), .B(_20589__bF_buf4), .C(_21294_), .Y(_21295_) );
	NOR2X1 NOR2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_21293_), .B(_21295_), .Y(_21296_) );
	NAND3X1 NAND3X1_3901 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_20_), .B(bLoc_frameOut_4_bF_buf2), .C(_20595__bF_buf4), .Y(_21297_) );
	OAI21X1 OAI21X1_4743 ( .gnd(gnd), .vdd(vdd), .A(_18520_), .B(_20594__bF_buf4), .C(_21297_), .Y(_21298_) );
	NAND3X1 NAND3X1_3902 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_20_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_21299_) );
	OAI21X1 OAI21X1_4744 ( .gnd(gnd), .vdd(vdd), .A(_18523_), .B(_20598__bF_buf4), .C(_21299_), .Y(_21300_) );
	NOR2X1 NOR2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_21298_), .B(_21300_), .Y(_21301_) );
	NAND2X1 NAND2X1_3681 ( .gnd(gnd), .vdd(vdd), .A(_21301_), .B(_21296_), .Y(_21302_) );
	NOR2X1 NOR2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_21302_), .B(_21292_), .Y(_21303_) );
	AOI22X1 AOI22X1_482 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_20_), .C(registers_r1_20_), .D(_20606__bF_buf4), .Y(_21304_) );
	AOI22X1 AOI22X1_483 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_20_), .C(registers_r5_20_), .D(_20611__bF_buf4), .Y(_21305_) );
	NAND3X1 NAND3X1_3903 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_20_), .B(_20607__bF_buf2), .C(_20574__bF_buf1), .Y(_21306_) );
	OAI21X1 OAI21X1_4745 ( .gnd(gnd), .vdd(vdd), .A(_18531_), .B(_20617__bF_buf4), .C(_21306_), .Y(_21307_) );
	AOI21X1 AOI21X1_3167 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_20_), .B(_20615__bF_buf4), .C(_21307_), .Y(_21308_) );
	NAND3X1 NAND3X1_3904 ( .gnd(gnd), .vdd(vdd), .A(_21304_), .B(_21305_), .C(_21308_), .Y(_21309_) );
	OAI22X1 OAI22X1_572 ( .gnd(gnd), .vdd(vdd), .A(_18537_), .B(_20622__bF_buf4), .C(_18536_), .D(_20621__bF_buf4), .Y(_21310_) );
	OAI22X1 OAI22X1_573 ( .gnd(gnd), .vdd(vdd), .A(_18539_), .B(_20626__bF_buf4), .C(_18540_), .D(_20624__bF_buf4), .Y(_21311_) );
	NOR2X1 NOR2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_21311_), .B(_21310_), .Y(_21312_) );
	OAI22X1 OAI22X1_574 ( .gnd(gnd), .vdd(vdd), .A(_18543_), .B(_20629__bF_buf4), .C(_18544_), .D(_20630__bF_buf4), .Y(_21313_) );
	OAI22X1 OAI22X1_575 ( .gnd(gnd), .vdd(vdd), .A(_18547_), .B(_20633__bF_buf4), .C(_18546_), .D(_20632__bF_buf4), .Y(_21314_) );
	NOR2X1 NOR2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_21313_), .B(_21314_), .Y(_21315_) );
	NAND2X1 NAND2X1_3682 ( .gnd(gnd), .vdd(vdd), .A(_21312_), .B(_21315_), .Y(_21316_) );
	NOR2X1 NOR2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_21309_), .B(_21316_), .Y(_21317_) );
	NAND2X1 NAND2X1_3683 ( .gnd(gnd), .vdd(vdd), .A(_21317_), .B(_21303_), .Y(readB_regOut_20_) );
	NAND3X1 NAND3X1_3905 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_21_), .B(_20559__bF_buf2), .C(_20557__bF_buf4), .Y(_21318_) );
	NAND3X1 NAND3X1_3906 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_21_), .B(_20562__bF_buf2), .C(_20557__bF_buf3), .Y(_21319_) );
	NAND2X1 NAND2X1_3684 ( .gnd(gnd), .vdd(vdd), .A(_21318_), .B(_21319_), .Y(_21320_) );
	OAI22X1 OAI22X1_576 ( .gnd(gnd), .vdd(vdd), .A(_18555_), .B(_20568__bF_buf3), .C(_18556_), .D(_20567__bF_buf3), .Y(_21321_) );
	NOR2X1 NOR2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_21320_), .B(_21321_), .Y(_21322_) );
	OAI22X1 OAI22X1_577 ( .gnd(gnd), .vdd(vdd), .A(_18559_), .B(_20576__bF_buf3), .C(_18560_), .D(_20575__bF_buf3), .Y(_21323_) );
	OAI22X1 OAI22X1_578 ( .gnd(gnd), .vdd(vdd), .A(_18562_), .B(_20581__bF_buf3), .C(_18563_), .D(_20580__bF_buf3), .Y(_21324_) );
	NOR2X1 NOR2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_21324_), .B(_21323_), .Y(_21325_) );
	NAND2X1 NAND2X1_3685 ( .gnd(gnd), .vdd(vdd), .A(_21322_), .B(_21325_), .Y(_21326_) );
	OAI22X1 OAI22X1_579 ( .gnd(gnd), .vdd(vdd), .A(_18568_), .B(_20586__bF_buf3), .C(_18567_), .D(_20585__bF_buf3), .Y(_21327_) );
	NAND3X1 NAND3X1_3907 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_21_), .B(_20588__bF_buf4), .C(_20590__bF_buf5), .Y(_21328_) );
	OAI21X1 OAI21X1_4746 ( .gnd(gnd), .vdd(vdd), .A(_18570_), .B(_20589__bF_buf3), .C(_21328_), .Y(_21329_) );
	NOR2X1 NOR2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_21327_), .B(_21329_), .Y(_21330_) );
	NAND3X1 NAND3X1_3908 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_21_), .B(bLoc_frameOut_4_bF_buf1), .C(_20595__bF_buf3), .Y(_21331_) );
	OAI21X1 OAI21X1_4747 ( .gnd(gnd), .vdd(vdd), .A(_18574_), .B(_20594__bF_buf3), .C(_21331_), .Y(_21332_) );
	NAND3X1 NAND3X1_3909 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_21_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_21333_) );
	OAI21X1 OAI21X1_4748 ( .gnd(gnd), .vdd(vdd), .A(_18577_), .B(_20598__bF_buf3), .C(_21333_), .Y(_21334_) );
	NOR2X1 NOR2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_21332_), .B(_21334_), .Y(_21335_) );
	NAND2X1 NAND2X1_3686 ( .gnd(gnd), .vdd(vdd), .A(_21335_), .B(_21330_), .Y(_21336_) );
	NOR2X1 NOR2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_21336_), .B(_21326_), .Y(_21337_) );
	AOI22X1 AOI22X1_484 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_21_), .C(registers_r1_21_), .D(_20606__bF_buf3), .Y(_21338_) );
	AOI22X1 AOI22X1_485 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_21_), .C(registers_r5_21_), .D(_20611__bF_buf3), .Y(_21339_) );
	NAND3X1 NAND3X1_3910 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_21_), .B(_20607__bF_buf1), .C(_20574__bF_buf7), .Y(_21340_) );
	OAI21X1 OAI21X1_4749 ( .gnd(gnd), .vdd(vdd), .A(_18585_), .B(_20617__bF_buf3), .C(_21340_), .Y(_21341_) );
	AOI21X1 AOI21X1_3168 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_21_), .B(_20615__bF_buf3), .C(_21341_), .Y(_21342_) );
	NAND3X1 NAND3X1_3911 ( .gnd(gnd), .vdd(vdd), .A(_21338_), .B(_21339_), .C(_21342_), .Y(_21343_) );
	OAI22X1 OAI22X1_580 ( .gnd(gnd), .vdd(vdd), .A(_18591_), .B(_20622__bF_buf3), .C(_18590_), .D(_20621__bF_buf3), .Y(_21344_) );
	OAI22X1 OAI22X1_581 ( .gnd(gnd), .vdd(vdd), .A(_18593_), .B(_20626__bF_buf3), .C(_18594_), .D(_20624__bF_buf3), .Y(_21345_) );
	NOR2X1 NOR2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_21345_), .B(_21344_), .Y(_21346_) );
	OAI22X1 OAI22X1_582 ( .gnd(gnd), .vdd(vdd), .A(_18597_), .B(_20629__bF_buf3), .C(_18598_), .D(_20630__bF_buf3), .Y(_21347_) );
	OAI22X1 OAI22X1_583 ( .gnd(gnd), .vdd(vdd), .A(_18601_), .B(_20633__bF_buf3), .C(_18600_), .D(_20632__bF_buf3), .Y(_21348_) );
	NOR2X1 NOR2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_21347_), .B(_21348_), .Y(_21349_) );
	NAND2X1 NAND2X1_3687 ( .gnd(gnd), .vdd(vdd), .A(_21346_), .B(_21349_), .Y(_21350_) );
	NOR2X1 NOR2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_21343_), .B(_21350_), .Y(_21351_) );
	NAND2X1 NAND2X1_3688 ( .gnd(gnd), .vdd(vdd), .A(_21351_), .B(_21337_), .Y(readB_regOut_21_) );
	NAND3X1 NAND3X1_3912 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_22_), .B(_20559__bF_buf1), .C(_20557__bF_buf2), .Y(_21352_) );
	NAND3X1 NAND3X1_3913 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_22_), .B(_20562__bF_buf1), .C(_20557__bF_buf1), .Y(_21353_) );
	NAND2X1 NAND2X1_3689 ( .gnd(gnd), .vdd(vdd), .A(_21352_), .B(_21353_), .Y(_21354_) );
	OAI22X1 OAI22X1_584 ( .gnd(gnd), .vdd(vdd), .A(_18609_), .B(_20568__bF_buf2), .C(_18610_), .D(_20567__bF_buf2), .Y(_21355_) );
	NOR2X1 NOR2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_21354_), .B(_21355_), .Y(_21356_) );
	OAI22X1 OAI22X1_585 ( .gnd(gnd), .vdd(vdd), .A(_18613_), .B(_20576__bF_buf2), .C(_18614_), .D(_20575__bF_buf2), .Y(_21357_) );
	OAI22X1 OAI22X1_586 ( .gnd(gnd), .vdd(vdd), .A(_18616_), .B(_20581__bF_buf2), .C(_18617_), .D(_20580__bF_buf2), .Y(_21358_) );
	NOR2X1 NOR2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_21358_), .B(_21357_), .Y(_21359_) );
	NAND2X1 NAND2X1_3690 ( .gnd(gnd), .vdd(vdd), .A(_21356_), .B(_21359_), .Y(_21360_) );
	OAI22X1 OAI22X1_587 ( .gnd(gnd), .vdd(vdd), .A(_18622_), .B(_20586__bF_buf2), .C(_18621_), .D(_20585__bF_buf2), .Y(_21361_) );
	NAND3X1 NAND3X1_3914 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_22_), .B(_20588__bF_buf3), .C(_20590__bF_buf3), .Y(_21362_) );
	OAI21X1 OAI21X1_4750 ( .gnd(gnd), .vdd(vdd), .A(_18624_), .B(_20589__bF_buf2), .C(_21362_), .Y(_21363_) );
	NOR2X1 NOR2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_21361_), .B(_21363_), .Y(_21364_) );
	NAND3X1 NAND3X1_3915 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_22_), .B(bLoc_frameOut_4_bF_buf0), .C(_20595__bF_buf2), .Y(_21365_) );
	OAI21X1 OAI21X1_4751 ( .gnd(gnd), .vdd(vdd), .A(_18628_), .B(_20594__bF_buf2), .C(_21365_), .Y(_21366_) );
	NAND3X1 NAND3X1_3916 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_22_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_21367_) );
	OAI21X1 OAI21X1_4752 ( .gnd(gnd), .vdd(vdd), .A(_18631_), .B(_20598__bF_buf2), .C(_21367_), .Y(_21368_) );
	NOR2X1 NOR2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_21366_), .B(_21368_), .Y(_21369_) );
	NAND2X1 NAND2X1_3691 ( .gnd(gnd), .vdd(vdd), .A(_21369_), .B(_21364_), .Y(_21370_) );
	NOR2X1 NOR2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_21370_), .B(_21360_), .Y(_21371_) );
	AOI22X1 AOI22X1_486 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf2), .B(registers_a2_22_), .C(registers_r1_22_), .D(_20606__bF_buf2), .Y(_21372_) );
	AOI22X1 AOI22X1_487 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf2), .B(registers_r4_22_), .C(registers_r5_22_), .D(_20611__bF_buf2), .Y(_21373_) );
	NAND3X1 NAND3X1_3917 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_22_), .B(_20607__bF_buf0), .C(_20574__bF_buf5), .Y(_21374_) );
	OAI21X1 OAI21X1_4753 ( .gnd(gnd), .vdd(vdd), .A(_18639_), .B(_20617__bF_buf2), .C(_21374_), .Y(_21375_) );
	AOI21X1 AOI21X1_3169 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_22_), .B(_20615__bF_buf2), .C(_21375_), .Y(_21376_) );
	NAND3X1 NAND3X1_3918 ( .gnd(gnd), .vdd(vdd), .A(_21372_), .B(_21373_), .C(_21376_), .Y(_21377_) );
	OAI22X1 OAI22X1_588 ( .gnd(gnd), .vdd(vdd), .A(_18645_), .B(_20622__bF_buf2), .C(_18644_), .D(_20621__bF_buf2), .Y(_21378_) );
	OAI22X1 OAI22X1_589 ( .gnd(gnd), .vdd(vdd), .A(_18647_), .B(_20626__bF_buf2), .C(_18648_), .D(_20624__bF_buf2), .Y(_21379_) );
	NOR2X1 NOR2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_21379_), .B(_21378_), .Y(_21380_) );
	OAI22X1 OAI22X1_590 ( .gnd(gnd), .vdd(vdd), .A(_18651_), .B(_20629__bF_buf2), .C(_18652_), .D(_20630__bF_buf2), .Y(_21381_) );
	OAI22X1 OAI22X1_591 ( .gnd(gnd), .vdd(vdd), .A(_18655_), .B(_20633__bF_buf2), .C(_18654_), .D(_20632__bF_buf2), .Y(_21382_) );
	NOR2X1 NOR2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_21381_), .B(_21382_), .Y(_21383_) );
	NAND2X1 NAND2X1_3692 ( .gnd(gnd), .vdd(vdd), .A(_21380_), .B(_21383_), .Y(_21384_) );
	NOR2X1 NOR2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_21377_), .B(_21384_), .Y(_21385_) );
	NAND2X1 NAND2X1_3693 ( .gnd(gnd), .vdd(vdd), .A(_21385_), .B(_21371_), .Y(readB_regOut_22_) );
	NAND3X1 NAND3X1_3919 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_23_), .B(_20559__bF_buf0), .C(_20557__bF_buf0), .Y(_21386_) );
	NAND3X1 NAND3X1_3920 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_23_), .B(_20562__bF_buf0), .C(_20557__bF_buf7), .Y(_21387_) );
	NAND2X1 NAND2X1_3694 ( .gnd(gnd), .vdd(vdd), .A(_21386_), .B(_21387_), .Y(_21388_) );
	OAI22X1 OAI22X1_592 ( .gnd(gnd), .vdd(vdd), .A(_18663_), .B(_20568__bF_buf1), .C(_18664_), .D(_20567__bF_buf1), .Y(_21389_) );
	NOR2X1 NOR2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_21388_), .B(_21389_), .Y(_21390_) );
	OAI22X1 OAI22X1_593 ( .gnd(gnd), .vdd(vdd), .A(_18667_), .B(_20576__bF_buf1), .C(_18668_), .D(_20575__bF_buf1), .Y(_21391_) );
	OAI22X1 OAI22X1_594 ( .gnd(gnd), .vdd(vdd), .A(_18670_), .B(_20581__bF_buf1), .C(_18671_), .D(_20580__bF_buf1), .Y(_21392_) );
	NOR2X1 NOR2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_21392_), .B(_21391_), .Y(_21393_) );
	NAND2X1 NAND2X1_3695 ( .gnd(gnd), .vdd(vdd), .A(_21390_), .B(_21393_), .Y(_21394_) );
	OAI22X1 OAI22X1_595 ( .gnd(gnd), .vdd(vdd), .A(_18676_), .B(_20586__bF_buf1), .C(_18675_), .D(_20585__bF_buf1), .Y(_21395_) );
	NAND3X1 NAND3X1_3921 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_23_), .B(_20588__bF_buf2), .C(_20590__bF_buf1), .Y(_21396_) );
	OAI21X1 OAI21X1_4754 ( .gnd(gnd), .vdd(vdd), .A(_18678_), .B(_20589__bF_buf1), .C(_21396_), .Y(_21397_) );
	NOR2X1 NOR2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_21395_), .B(_21397_), .Y(_21398_) );
	NAND3X1 NAND3X1_3922 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_23_), .B(bLoc_frameOut_4_bF_buf6), .C(_20595__bF_buf1), .Y(_21399_) );
	OAI21X1 OAI21X1_4755 ( .gnd(gnd), .vdd(vdd), .A(_18682_), .B(_20594__bF_buf1), .C(_21399_), .Y(_21400_) );
	NAND3X1 NAND3X1_3923 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_23_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_21401_) );
	OAI21X1 OAI21X1_4756 ( .gnd(gnd), .vdd(vdd), .A(_18685_), .B(_20598__bF_buf1), .C(_21401_), .Y(_21402_) );
	NOR2X1 NOR2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_21400_), .B(_21402_), .Y(_21403_) );
	NAND2X1 NAND2X1_3696 ( .gnd(gnd), .vdd(vdd), .A(_21403_), .B(_21398_), .Y(_21404_) );
	NOR2X1 NOR2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_21404_), .B(_21394_), .Y(_21405_) );
	AOI22X1 AOI22X1_488 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf1), .B(registers_a2_23_), .C(registers_r1_23_), .D(_20606__bF_buf1), .Y(_21406_) );
	AOI22X1 AOI22X1_489 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf1), .B(registers_r4_23_), .C(registers_r5_23_), .D(_20611__bF_buf1), .Y(_21407_) );
	NAND3X1 NAND3X1_3924 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_23_), .B(_20607__bF_buf4), .C(_20574__bF_buf3), .Y(_21408_) );
	OAI21X1 OAI21X1_4757 ( .gnd(gnd), .vdd(vdd), .A(_18693_), .B(_20617__bF_buf1), .C(_21408_), .Y(_21409_) );
	AOI21X1 AOI21X1_3170 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_23_), .B(_20615__bF_buf1), .C(_21409_), .Y(_21410_) );
	NAND3X1 NAND3X1_3925 ( .gnd(gnd), .vdd(vdd), .A(_21406_), .B(_21407_), .C(_21410_), .Y(_21411_) );
	OAI22X1 OAI22X1_596 ( .gnd(gnd), .vdd(vdd), .A(_18699_), .B(_20622__bF_buf1), .C(_18698_), .D(_20621__bF_buf1), .Y(_21412_) );
	OAI22X1 OAI22X1_597 ( .gnd(gnd), .vdd(vdd), .A(_18701_), .B(_20626__bF_buf1), .C(_18702_), .D(_20624__bF_buf1), .Y(_21413_) );
	NOR2X1 NOR2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_21413_), .B(_21412_), .Y(_21414_) );
	OAI22X1 OAI22X1_598 ( .gnd(gnd), .vdd(vdd), .A(_18705_), .B(_20629__bF_buf1), .C(_18706_), .D(_20630__bF_buf1), .Y(_21415_) );
	OAI22X1 OAI22X1_599 ( .gnd(gnd), .vdd(vdd), .A(_18709_), .B(_20633__bF_buf1), .C(_18708_), .D(_20632__bF_buf1), .Y(_21416_) );
	NOR2X1 NOR2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_21415_), .B(_21416_), .Y(_21417_) );
	NAND2X1 NAND2X1_3697 ( .gnd(gnd), .vdd(vdd), .A(_21414_), .B(_21417_), .Y(_21418_) );
	NOR2X1 NOR2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_21411_), .B(_21418_), .Y(_21419_) );
	NAND2X1 NAND2X1_3698 ( .gnd(gnd), .vdd(vdd), .A(_21419_), .B(_21405_), .Y(readB_regOut_23_) );
	NAND3X1 NAND3X1_3926 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_24_), .B(_20559__bF_buf5), .C(_20557__bF_buf6), .Y(_21420_) );
	NAND3X1 NAND3X1_3927 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_24_), .B(_20562__bF_buf5), .C(_20557__bF_buf5), .Y(_21421_) );
	NAND2X1 NAND2X1_3699 ( .gnd(gnd), .vdd(vdd), .A(_21420_), .B(_21421_), .Y(_21422_) );
	OAI22X1 OAI22X1_600 ( .gnd(gnd), .vdd(vdd), .A(_18717_), .B(_20568__bF_buf0), .C(_18718_), .D(_20567__bF_buf0), .Y(_21423_) );
	NOR2X1 NOR2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_21422_), .B(_21423_), .Y(_21424_) );
	OAI22X1 OAI22X1_601 ( .gnd(gnd), .vdd(vdd), .A(_18721_), .B(_20576__bF_buf0), .C(_18722_), .D(_20575__bF_buf0), .Y(_21425_) );
	OAI22X1 OAI22X1_602 ( .gnd(gnd), .vdd(vdd), .A(_18724_), .B(_20581__bF_buf0), .C(_18725_), .D(_20580__bF_buf0), .Y(_21426_) );
	NOR2X1 NOR2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_21426_), .B(_21425_), .Y(_21427_) );
	NAND2X1 NAND2X1_3700 ( .gnd(gnd), .vdd(vdd), .A(_21424_), .B(_21427_), .Y(_21428_) );
	OAI22X1 OAI22X1_603 ( .gnd(gnd), .vdd(vdd), .A(_18730_), .B(_20586__bF_buf0), .C(_18729_), .D(_20585__bF_buf0), .Y(_21429_) );
	NAND3X1 NAND3X1_3928 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_24_), .B(_20588__bF_buf1), .C(_20590__bF_buf7), .Y(_21430_) );
	OAI21X1 OAI21X1_4758 ( .gnd(gnd), .vdd(vdd), .A(_18732_), .B(_20589__bF_buf0), .C(_21430_), .Y(_21431_) );
	NOR2X1 NOR2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_21429_), .B(_21431_), .Y(_21432_) );
	NAND3X1 NAND3X1_3929 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_24_), .B(bLoc_frameOut_4_bF_buf5), .C(_20595__bF_buf0), .Y(_21433_) );
	OAI21X1 OAI21X1_4759 ( .gnd(gnd), .vdd(vdd), .A(_18736_), .B(_20594__bF_buf0), .C(_21433_), .Y(_21434_) );
	NAND3X1 NAND3X1_3930 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_24_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_21435_) );
	OAI21X1 OAI21X1_4760 ( .gnd(gnd), .vdd(vdd), .A(_18739_), .B(_20598__bF_buf0), .C(_21435_), .Y(_21436_) );
	NOR2X1 NOR2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_21434_), .B(_21436_), .Y(_21437_) );
	NAND2X1 NAND2X1_3701 ( .gnd(gnd), .vdd(vdd), .A(_21437_), .B(_21432_), .Y(_21438_) );
	NOR2X1 NOR2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_21438_), .B(_21428_), .Y(_21439_) );
	AOI22X1 AOI22X1_490 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf0), .B(registers_a2_24_), .C(registers_r1_24_), .D(_20606__bF_buf0), .Y(_21440_) );
	AOI22X1 AOI22X1_491 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf0), .B(registers_r4_24_), .C(registers_r5_24_), .D(_20611__bF_buf0), .Y(_21441_) );
	NAND3X1 NAND3X1_3931 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_24_), .B(_20607__bF_buf3), .C(_20574__bF_buf1), .Y(_21442_) );
	OAI21X1 OAI21X1_4761 ( .gnd(gnd), .vdd(vdd), .A(_18747_), .B(_20617__bF_buf0), .C(_21442_), .Y(_21443_) );
	AOI21X1 AOI21X1_3171 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_24_), .B(_20615__bF_buf0), .C(_21443_), .Y(_21444_) );
	NAND3X1 NAND3X1_3932 ( .gnd(gnd), .vdd(vdd), .A(_21440_), .B(_21441_), .C(_21444_), .Y(_21445_) );
	OAI22X1 OAI22X1_604 ( .gnd(gnd), .vdd(vdd), .A(_18753_), .B(_20622__bF_buf0), .C(_18752_), .D(_20621__bF_buf0), .Y(_21446_) );
	OAI22X1 OAI22X1_605 ( .gnd(gnd), .vdd(vdd), .A(_18755_), .B(_20626__bF_buf0), .C(_18756_), .D(_20624__bF_buf0), .Y(_21447_) );
	NOR2X1 NOR2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_21447_), .B(_21446_), .Y(_21448_) );
	OAI22X1 OAI22X1_606 ( .gnd(gnd), .vdd(vdd), .A(_18759_), .B(_20629__bF_buf0), .C(_18760_), .D(_20630__bF_buf0), .Y(_21449_) );
	OAI22X1 OAI22X1_607 ( .gnd(gnd), .vdd(vdd), .A(_18763_), .B(_20633__bF_buf0), .C(_18762_), .D(_20632__bF_buf0), .Y(_21450_) );
	NOR2X1 NOR2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_21449_), .B(_21450_), .Y(_21451_) );
	NAND2X1 NAND2X1_3702 ( .gnd(gnd), .vdd(vdd), .A(_21448_), .B(_21451_), .Y(_21452_) );
	NOR2X1 NOR2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_21445_), .B(_21452_), .Y(_21453_) );
	NAND2X1 NAND2X1_3703 ( .gnd(gnd), .vdd(vdd), .A(_21453_), .B(_21439_), .Y(readB_regOut_24_) );
	NAND3X1 NAND3X1_3933 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_25_), .B(_20559__bF_buf4), .C(_20557__bF_buf4), .Y(_21454_) );
	NAND3X1 NAND3X1_3934 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_25_), .B(_20562__bF_buf4), .C(_20557__bF_buf3), .Y(_21455_) );
	NAND2X1 NAND2X1_3704 ( .gnd(gnd), .vdd(vdd), .A(_21454_), .B(_21455_), .Y(_21456_) );
	OAI22X1 OAI22X1_608 ( .gnd(gnd), .vdd(vdd), .A(_18771_), .B(_20568__bF_buf4), .C(_18772_), .D(_20567__bF_buf4), .Y(_21457_) );
	NOR2X1 NOR2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_21456_), .B(_21457_), .Y(_21458_) );
	OAI22X1 OAI22X1_609 ( .gnd(gnd), .vdd(vdd), .A(_18775_), .B(_20576__bF_buf4), .C(_18776_), .D(_20575__bF_buf4), .Y(_21459_) );
	OAI22X1 OAI22X1_610 ( .gnd(gnd), .vdd(vdd), .A(_18778_), .B(_20581__bF_buf4), .C(_18779_), .D(_20580__bF_buf4), .Y(_21460_) );
	NOR2X1 NOR2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_21460_), .B(_21459_), .Y(_21461_) );
	NAND2X1 NAND2X1_3705 ( .gnd(gnd), .vdd(vdd), .A(_21458_), .B(_21461_), .Y(_21462_) );
	OAI22X1 OAI22X1_611 ( .gnd(gnd), .vdd(vdd), .A(_18784_), .B(_20586__bF_buf4), .C(_18783_), .D(_20585__bF_buf4), .Y(_21463_) );
	NAND3X1 NAND3X1_3935 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_25_), .B(_20588__bF_buf0), .C(_20590__bF_buf5), .Y(_21464_) );
	OAI21X1 OAI21X1_4762 ( .gnd(gnd), .vdd(vdd), .A(_18786_), .B(_20589__bF_buf4), .C(_21464_), .Y(_21465_) );
	NOR2X1 NOR2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_21463_), .B(_21465_), .Y(_21466_) );
	NAND3X1 NAND3X1_3936 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_25_), .B(bLoc_frameOut_4_bF_buf4), .C(_20595__bF_buf4), .Y(_21467_) );
	OAI21X1 OAI21X1_4763 ( .gnd(gnd), .vdd(vdd), .A(_18790_), .B(_20594__bF_buf4), .C(_21467_), .Y(_21468_) );
	NAND3X1 NAND3X1_3937 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_25_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_21469_) );
	OAI21X1 OAI21X1_4764 ( .gnd(gnd), .vdd(vdd), .A(_18793_), .B(_20598__bF_buf4), .C(_21469_), .Y(_21470_) );
	NOR2X1 NOR2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_21468_), .B(_21470_), .Y(_21471_) );
	NAND2X1 NAND2X1_3706 ( .gnd(gnd), .vdd(vdd), .A(_21471_), .B(_21466_), .Y(_21472_) );
	NOR2X1 NOR2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_21472_), .B(_21462_), .Y(_21473_) );
	AOI22X1 AOI22X1_492 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_25_), .C(registers_r1_25_), .D(_20606__bF_buf4), .Y(_21474_) );
	AOI22X1 AOI22X1_493 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_25_), .C(registers_r5_25_), .D(_20611__bF_buf4), .Y(_21475_) );
	NAND3X1 NAND3X1_3938 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_25_), .B(_20607__bF_buf2), .C(_20574__bF_buf7), .Y(_21476_) );
	OAI21X1 OAI21X1_4765 ( .gnd(gnd), .vdd(vdd), .A(_18801_), .B(_20617__bF_buf4), .C(_21476_), .Y(_21477_) );
	AOI21X1 AOI21X1_3172 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_25_), .B(_20615__bF_buf4), .C(_21477_), .Y(_21478_) );
	NAND3X1 NAND3X1_3939 ( .gnd(gnd), .vdd(vdd), .A(_21474_), .B(_21475_), .C(_21478_), .Y(_21479_) );
	OAI22X1 OAI22X1_612 ( .gnd(gnd), .vdd(vdd), .A(_18807_), .B(_20622__bF_buf4), .C(_18806_), .D(_20621__bF_buf4), .Y(_21480_) );
	OAI22X1 OAI22X1_613 ( .gnd(gnd), .vdd(vdd), .A(_18809_), .B(_20626__bF_buf4), .C(_18810_), .D(_20624__bF_buf4), .Y(_21481_) );
	NOR2X1 NOR2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_21481_), .B(_21480_), .Y(_21482_) );
	OAI22X1 OAI22X1_614 ( .gnd(gnd), .vdd(vdd), .A(_18813_), .B(_20629__bF_buf4), .C(_18814_), .D(_20630__bF_buf4), .Y(_21483_) );
	OAI22X1 OAI22X1_615 ( .gnd(gnd), .vdd(vdd), .A(_18817_), .B(_20633__bF_buf4), .C(_18816_), .D(_20632__bF_buf4), .Y(_21484_) );
	NOR2X1 NOR2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_21483_), .B(_21484_), .Y(_21485_) );
	NAND2X1 NAND2X1_3707 ( .gnd(gnd), .vdd(vdd), .A(_21482_), .B(_21485_), .Y(_21486_) );
	NOR2X1 NOR2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_21479_), .B(_21486_), .Y(_21487_) );
	NAND2X1 NAND2X1_3708 ( .gnd(gnd), .vdd(vdd), .A(_21487_), .B(_21473_), .Y(readB_regOut_25_) );
	NAND3X1 NAND3X1_3940 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_26_), .B(_20559__bF_buf3), .C(_20557__bF_buf2), .Y(_21488_) );
	NAND3X1 NAND3X1_3941 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_26_), .B(_20562__bF_buf3), .C(_20557__bF_buf1), .Y(_21489_) );
	NAND2X1 NAND2X1_3709 ( .gnd(gnd), .vdd(vdd), .A(_21488_), .B(_21489_), .Y(_21490_) );
	OAI22X1 OAI22X1_616 ( .gnd(gnd), .vdd(vdd), .A(_18825_), .B(_20568__bF_buf3), .C(_18826_), .D(_20567__bF_buf3), .Y(_21491_) );
	NOR2X1 NOR2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_21490_), .B(_21491_), .Y(_21492_) );
	OAI22X1 OAI22X1_617 ( .gnd(gnd), .vdd(vdd), .A(_18829_), .B(_20576__bF_buf3), .C(_18830_), .D(_20575__bF_buf3), .Y(_21493_) );
	OAI22X1 OAI22X1_618 ( .gnd(gnd), .vdd(vdd), .A(_18832_), .B(_20581__bF_buf3), .C(_18833_), .D(_20580__bF_buf3), .Y(_21494_) );
	NOR2X1 NOR2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_21494_), .B(_21493_), .Y(_21495_) );
	NAND2X1 NAND2X1_3710 ( .gnd(gnd), .vdd(vdd), .A(_21492_), .B(_21495_), .Y(_21496_) );
	OAI22X1 OAI22X1_619 ( .gnd(gnd), .vdd(vdd), .A(_18838_), .B(_20586__bF_buf3), .C(_18837_), .D(_20585__bF_buf3), .Y(_21497_) );
	NAND3X1 NAND3X1_3942 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_26_), .B(_20588__bF_buf5), .C(_20590__bF_buf3), .Y(_21498_) );
	OAI21X1 OAI21X1_4766 ( .gnd(gnd), .vdd(vdd), .A(_18840_), .B(_20589__bF_buf3), .C(_21498_), .Y(_21499_) );
	NOR2X1 NOR2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_21497_), .B(_21499_), .Y(_21500_) );
	NAND3X1 NAND3X1_3943 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_26_), .B(bLoc_frameOut_4_bF_buf3), .C(_20595__bF_buf3), .Y(_21501_) );
	OAI21X1 OAI21X1_4767 ( .gnd(gnd), .vdd(vdd), .A(_18844_), .B(_20594__bF_buf3), .C(_21501_), .Y(_21502_) );
	NAND3X1 NAND3X1_3944 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_26_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_21503_) );
	OAI21X1 OAI21X1_4768 ( .gnd(gnd), .vdd(vdd), .A(_18847_), .B(_20598__bF_buf3), .C(_21503_), .Y(_21504_) );
	NOR2X1 NOR2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_21502_), .B(_21504_), .Y(_21505_) );
	NAND2X1 NAND2X1_3711 ( .gnd(gnd), .vdd(vdd), .A(_21505_), .B(_21500_), .Y(_21506_) );
	NOR2X1 NOR2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_21506_), .B(_21496_), .Y(_21507_) );
	AOI22X1 AOI22X1_494 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_26_), .C(registers_r1_26_), .D(_20606__bF_buf3), .Y(_21508_) );
	AOI22X1 AOI22X1_495 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_26_), .C(registers_r5_26_), .D(_20611__bF_buf3), .Y(_21509_) );
	NAND3X1 NAND3X1_3945 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_26_), .B(_20607__bF_buf1), .C(_20574__bF_buf5), .Y(_21510_) );
	OAI21X1 OAI21X1_4769 ( .gnd(gnd), .vdd(vdd), .A(_18855_), .B(_20617__bF_buf3), .C(_21510_), .Y(_21511_) );
	AOI21X1 AOI21X1_3173 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_26_), .B(_20615__bF_buf3), .C(_21511_), .Y(_21512_) );
	NAND3X1 NAND3X1_3946 ( .gnd(gnd), .vdd(vdd), .A(_21508_), .B(_21509_), .C(_21512_), .Y(_21513_) );
	OAI22X1 OAI22X1_620 ( .gnd(gnd), .vdd(vdd), .A(_18861_), .B(_20622__bF_buf3), .C(_18860_), .D(_20621__bF_buf3), .Y(_21514_) );
	OAI22X1 OAI22X1_621 ( .gnd(gnd), .vdd(vdd), .A(_18863_), .B(_20626__bF_buf3), .C(_18864_), .D(_20624__bF_buf3), .Y(_21515_) );
	NOR2X1 NOR2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_21515_), .B(_21514_), .Y(_21516_) );
	OAI22X1 OAI22X1_622 ( .gnd(gnd), .vdd(vdd), .A(_18867_), .B(_20629__bF_buf3), .C(_18868_), .D(_20630__bF_buf3), .Y(_21517_) );
	OAI22X1 OAI22X1_623 ( .gnd(gnd), .vdd(vdd), .A(_18871_), .B(_20633__bF_buf3), .C(_18870_), .D(_20632__bF_buf3), .Y(_21518_) );
	NOR2X1 NOR2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_21517_), .B(_21518_), .Y(_21519_) );
	NAND2X1 NAND2X1_3712 ( .gnd(gnd), .vdd(vdd), .A(_21516_), .B(_21519_), .Y(_21520_) );
	NOR2X1 NOR2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_21513_), .B(_21520_), .Y(_21521_) );
	NAND2X1 NAND2X1_3713 ( .gnd(gnd), .vdd(vdd), .A(_21521_), .B(_21507_), .Y(readB_regOut_26_) );
	NAND3X1 NAND3X1_3947 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_27_), .B(_20559__bF_buf2), .C(_20557__bF_buf0), .Y(_21522_) );
	NAND3X1 NAND3X1_3948 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_27_), .B(_20562__bF_buf2), .C(_20557__bF_buf7), .Y(_21523_) );
	NAND2X1 NAND2X1_3714 ( .gnd(gnd), .vdd(vdd), .A(_21522_), .B(_21523_), .Y(_21524_) );
	OAI22X1 OAI22X1_624 ( .gnd(gnd), .vdd(vdd), .A(_18879_), .B(_20568__bF_buf2), .C(_18880_), .D(_20567__bF_buf2), .Y(_21525_) );
	NOR2X1 NOR2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_21524_), .B(_21525_), .Y(_21526_) );
	OAI22X1 OAI22X1_625 ( .gnd(gnd), .vdd(vdd), .A(_18883_), .B(_20576__bF_buf2), .C(_18884_), .D(_20575__bF_buf2), .Y(_21527_) );
	OAI22X1 OAI22X1_626 ( .gnd(gnd), .vdd(vdd), .A(_18886_), .B(_20581__bF_buf2), .C(_18887_), .D(_20580__bF_buf2), .Y(_21528_) );
	NOR2X1 NOR2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_21528_), .B(_21527_), .Y(_21529_) );
	NAND2X1 NAND2X1_3715 ( .gnd(gnd), .vdd(vdd), .A(_21526_), .B(_21529_), .Y(_21530_) );
	OAI22X1 OAI22X1_627 ( .gnd(gnd), .vdd(vdd), .A(_18892_), .B(_20586__bF_buf2), .C(_18891_), .D(_20585__bF_buf2), .Y(_21531_) );
	NAND3X1 NAND3X1_3949 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_27_), .B(_20588__bF_buf4), .C(_20590__bF_buf1), .Y(_21532_) );
	OAI21X1 OAI21X1_4770 ( .gnd(gnd), .vdd(vdd), .A(_18894_), .B(_20589__bF_buf2), .C(_21532_), .Y(_21533_) );
	NOR2X1 NOR2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_21531_), .B(_21533_), .Y(_21534_) );
	NAND3X1 NAND3X1_3950 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_27_), .B(bLoc_frameOut_4_bF_buf2), .C(_20595__bF_buf2), .Y(_21535_) );
	OAI21X1 OAI21X1_4771 ( .gnd(gnd), .vdd(vdd), .A(_18898_), .B(_20594__bF_buf2), .C(_21535_), .Y(_21536_) );
	NAND3X1 NAND3X1_3951 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_27_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_21537_) );
	OAI21X1 OAI21X1_4772 ( .gnd(gnd), .vdd(vdd), .A(_18901_), .B(_20598__bF_buf2), .C(_21537_), .Y(_21538_) );
	NOR2X1 NOR2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_21536_), .B(_21538_), .Y(_21539_) );
	NAND2X1 NAND2X1_3716 ( .gnd(gnd), .vdd(vdd), .A(_21539_), .B(_21534_), .Y(_21540_) );
	NOR2X1 NOR2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_21540_), .B(_21530_), .Y(_21541_) );
	AOI22X1 AOI22X1_496 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf2), .B(registers_a2_27_), .C(registers_r1_27_), .D(_20606__bF_buf2), .Y(_21542_) );
	AOI22X1 AOI22X1_497 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf2), .B(registers_r4_27_), .C(registers_r5_27_), .D(_20611__bF_buf2), .Y(_21543_) );
	NAND3X1 NAND3X1_3952 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_27_), .B(_20607__bF_buf0), .C(_20574__bF_buf3), .Y(_21544_) );
	OAI21X1 OAI21X1_4773 ( .gnd(gnd), .vdd(vdd), .A(_18909_), .B(_20617__bF_buf2), .C(_21544_), .Y(_21545_) );
	AOI21X1 AOI21X1_3174 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_27_), .B(_20615__bF_buf2), .C(_21545_), .Y(_21546_) );
	NAND3X1 NAND3X1_3953 ( .gnd(gnd), .vdd(vdd), .A(_21542_), .B(_21543_), .C(_21546_), .Y(_21547_) );
	OAI22X1 OAI22X1_628 ( .gnd(gnd), .vdd(vdd), .A(_18915_), .B(_20622__bF_buf2), .C(_18914_), .D(_20621__bF_buf2), .Y(_21548_) );
	OAI22X1 OAI22X1_629 ( .gnd(gnd), .vdd(vdd), .A(_18917_), .B(_20626__bF_buf2), .C(_18918_), .D(_20624__bF_buf2), .Y(_21549_) );
	NOR2X1 NOR2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_21549_), .B(_21548_), .Y(_21550_) );
	OAI22X1 OAI22X1_630 ( .gnd(gnd), .vdd(vdd), .A(_18921_), .B(_20629__bF_buf2), .C(_18922_), .D(_20630__bF_buf2), .Y(_21551_) );
	OAI22X1 OAI22X1_631 ( .gnd(gnd), .vdd(vdd), .A(_18925_), .B(_20633__bF_buf2), .C(_18924_), .D(_20632__bF_buf2), .Y(_21552_) );
	NOR2X1 NOR2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_21551_), .B(_21552_), .Y(_21553_) );
	NAND2X1 NAND2X1_3717 ( .gnd(gnd), .vdd(vdd), .A(_21550_), .B(_21553_), .Y(_21554_) );
	NOR2X1 NOR2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_21547_), .B(_21554_), .Y(_21555_) );
	NAND2X1 NAND2X1_3718 ( .gnd(gnd), .vdd(vdd), .A(_21555_), .B(_21541_), .Y(readB_regOut_27_) );
	NAND3X1 NAND3X1_3954 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_28_), .B(_20559__bF_buf1), .C(_20557__bF_buf6), .Y(_21556_) );
	NAND3X1 NAND3X1_3955 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_28_), .B(_20562__bF_buf1), .C(_20557__bF_buf5), .Y(_21557_) );
	NAND2X1 NAND2X1_3719 ( .gnd(gnd), .vdd(vdd), .A(_21556_), .B(_21557_), .Y(_21558_) );
	OAI22X1 OAI22X1_632 ( .gnd(gnd), .vdd(vdd), .A(_18933_), .B(_20568__bF_buf1), .C(_18934_), .D(_20567__bF_buf1), .Y(_21559_) );
	NOR2X1 NOR2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_21558_), .B(_21559_), .Y(_21560_) );
	OAI22X1 OAI22X1_633 ( .gnd(gnd), .vdd(vdd), .A(_18937_), .B(_20576__bF_buf1), .C(_18938_), .D(_20575__bF_buf1), .Y(_21561_) );
	OAI22X1 OAI22X1_634 ( .gnd(gnd), .vdd(vdd), .A(_18940_), .B(_20581__bF_buf1), .C(_18941_), .D(_20580__bF_buf1), .Y(_21562_) );
	NOR2X1 NOR2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_21562_), .B(_21561_), .Y(_21563_) );
	NAND2X1 NAND2X1_3720 ( .gnd(gnd), .vdd(vdd), .A(_21560_), .B(_21563_), .Y(_21564_) );
	OAI22X1 OAI22X1_635 ( .gnd(gnd), .vdd(vdd), .A(_18946_), .B(_20586__bF_buf1), .C(_18945_), .D(_20585__bF_buf1), .Y(_21565_) );
	NAND3X1 NAND3X1_3956 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_28_), .B(_20588__bF_buf3), .C(_20590__bF_buf7), .Y(_21566_) );
	OAI21X1 OAI21X1_4774 ( .gnd(gnd), .vdd(vdd), .A(_18948_), .B(_20589__bF_buf1), .C(_21566_), .Y(_21567_) );
	NOR2X1 NOR2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_21565_), .B(_21567_), .Y(_21568_) );
	NAND3X1 NAND3X1_3957 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_28_), .B(bLoc_frameOut_4_bF_buf1), .C(_20595__bF_buf1), .Y(_21569_) );
	OAI21X1 OAI21X1_4775 ( .gnd(gnd), .vdd(vdd), .A(_18952_), .B(_20594__bF_buf1), .C(_21569_), .Y(_21570_) );
	NAND3X1 NAND3X1_3958 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_28_), .B(_20574__bF_buf2), .C(_20590__bF_buf6), .Y(_21571_) );
	OAI21X1 OAI21X1_4776 ( .gnd(gnd), .vdd(vdd), .A(_18955_), .B(_20598__bF_buf1), .C(_21571_), .Y(_21572_) );
	NOR2X1 NOR2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_21570_), .B(_21572_), .Y(_21573_) );
	NAND2X1 NAND2X1_3721 ( .gnd(gnd), .vdd(vdd), .A(_21573_), .B(_21568_), .Y(_21574_) );
	NOR2X1 NOR2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_21574_), .B(_21564_), .Y(_21575_) );
	AOI22X1 AOI22X1_498 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf1), .B(registers_a2_28_), .C(registers_r1_28_), .D(_20606__bF_buf1), .Y(_21576_) );
	AOI22X1 AOI22X1_499 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf1), .B(registers_r4_28_), .C(registers_r5_28_), .D(_20611__bF_buf1), .Y(_21577_) );
	NAND3X1 NAND3X1_3959 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_28_), .B(_20607__bF_buf4), .C(_20574__bF_buf1), .Y(_21578_) );
	OAI21X1 OAI21X1_4777 ( .gnd(gnd), .vdd(vdd), .A(_18963_), .B(_20617__bF_buf1), .C(_21578_), .Y(_21579_) );
	AOI21X1 AOI21X1_3175 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_28_), .B(_20615__bF_buf1), .C(_21579_), .Y(_21580_) );
	NAND3X1 NAND3X1_3960 ( .gnd(gnd), .vdd(vdd), .A(_21576_), .B(_21577_), .C(_21580_), .Y(_21581_) );
	OAI22X1 OAI22X1_636 ( .gnd(gnd), .vdd(vdd), .A(_18969_), .B(_20622__bF_buf1), .C(_18968_), .D(_20621__bF_buf1), .Y(_21582_) );
	OAI22X1 OAI22X1_637 ( .gnd(gnd), .vdd(vdd), .A(_18971_), .B(_20626__bF_buf1), .C(_18972_), .D(_20624__bF_buf1), .Y(_21583_) );
	NOR2X1 NOR2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_21583_), .B(_21582_), .Y(_21584_) );
	OAI22X1 OAI22X1_638 ( .gnd(gnd), .vdd(vdd), .A(_18975_), .B(_20629__bF_buf1), .C(_18976_), .D(_20630__bF_buf1), .Y(_21585_) );
	OAI22X1 OAI22X1_639 ( .gnd(gnd), .vdd(vdd), .A(_18979_), .B(_20633__bF_buf1), .C(_18978_), .D(_20632__bF_buf1), .Y(_21586_) );
	NOR2X1 NOR2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_21585_), .B(_21586_), .Y(_21587_) );
	NAND2X1 NAND2X1_3722 ( .gnd(gnd), .vdd(vdd), .A(_21584_), .B(_21587_), .Y(_21588_) );
	NOR2X1 NOR2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_21581_), .B(_21588_), .Y(_21589_) );
	NAND2X1 NAND2X1_3723 ( .gnd(gnd), .vdd(vdd), .A(_21589_), .B(_21575_), .Y(readB_regOut_28_) );
	NAND3X1 NAND3X1_3961 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_29_), .B(_20559__bF_buf0), .C(_20557__bF_buf4), .Y(_21590_) );
	NAND3X1 NAND3X1_3962 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_29_), .B(_20562__bF_buf0), .C(_20557__bF_buf3), .Y(_21591_) );
	NAND2X1 NAND2X1_3724 ( .gnd(gnd), .vdd(vdd), .A(_21590_), .B(_21591_), .Y(_21592_) );
	OAI22X1 OAI22X1_640 ( .gnd(gnd), .vdd(vdd), .A(_18987_), .B(_20568__bF_buf0), .C(_18988_), .D(_20567__bF_buf0), .Y(_21593_) );
	NOR2X1 NOR2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_21592_), .B(_21593_), .Y(_21594_) );
	OAI22X1 OAI22X1_641 ( .gnd(gnd), .vdd(vdd), .A(_18991_), .B(_20576__bF_buf0), .C(_18992_), .D(_20575__bF_buf0), .Y(_21595_) );
	OAI22X1 OAI22X1_642 ( .gnd(gnd), .vdd(vdd), .A(_18994_), .B(_20581__bF_buf0), .C(_18995_), .D(_20580__bF_buf0), .Y(_21596_) );
	NOR2X1 NOR2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_21596_), .B(_21595_), .Y(_21597_) );
	NAND2X1 NAND2X1_3725 ( .gnd(gnd), .vdd(vdd), .A(_21594_), .B(_21597_), .Y(_21598_) );
	OAI22X1 OAI22X1_643 ( .gnd(gnd), .vdd(vdd), .A(_19000_), .B(_20586__bF_buf0), .C(_18999_), .D(_20585__bF_buf0), .Y(_21599_) );
	NAND3X1 NAND3X1_3963 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_29_), .B(_20588__bF_buf2), .C(_20590__bF_buf5), .Y(_21600_) );
	OAI21X1 OAI21X1_4778 ( .gnd(gnd), .vdd(vdd), .A(_19002_), .B(_20589__bF_buf0), .C(_21600_), .Y(_21601_) );
	NOR2X1 NOR2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_21599_), .B(_21601_), .Y(_21602_) );
	NAND3X1 NAND3X1_3964 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_29_), .B(bLoc_frameOut_4_bF_buf0), .C(_20595__bF_buf0), .Y(_21603_) );
	OAI21X1 OAI21X1_4779 ( .gnd(gnd), .vdd(vdd), .A(_19006_), .B(_20594__bF_buf0), .C(_21603_), .Y(_21604_) );
	NAND3X1 NAND3X1_3965 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_29_), .B(_20574__bF_buf0), .C(_20590__bF_buf4), .Y(_21605_) );
	OAI21X1 OAI21X1_4780 ( .gnd(gnd), .vdd(vdd), .A(_19009_), .B(_20598__bF_buf0), .C(_21605_), .Y(_21606_) );
	NOR2X1 NOR2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_21604_), .B(_21606_), .Y(_21607_) );
	NAND2X1 NAND2X1_3726 ( .gnd(gnd), .vdd(vdd), .A(_21607_), .B(_21602_), .Y(_21608_) );
	NOR2X1 NOR2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_21608_), .B(_21598_), .Y(_21609_) );
	AOI22X1 AOI22X1_500 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf0), .B(registers_a2_29_), .C(registers_r1_29_), .D(_20606__bF_buf0), .Y(_21610_) );
	AOI22X1 AOI22X1_501 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf0), .B(registers_r4_29_), .C(registers_r5_29_), .D(_20611__bF_buf0), .Y(_21611_) );
	NAND3X1 NAND3X1_3966 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_29_), .B(_20607__bF_buf3), .C(_20574__bF_buf7), .Y(_21612_) );
	OAI21X1 OAI21X1_4781 ( .gnd(gnd), .vdd(vdd), .A(_19017_), .B(_20617__bF_buf0), .C(_21612_), .Y(_21613_) );
	AOI21X1 AOI21X1_3176 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_29_), .B(_20615__bF_buf0), .C(_21613_), .Y(_21614_) );
	NAND3X1 NAND3X1_3967 ( .gnd(gnd), .vdd(vdd), .A(_21610_), .B(_21611_), .C(_21614_), .Y(_21615_) );
	OAI22X1 OAI22X1_644 ( .gnd(gnd), .vdd(vdd), .A(_19023_), .B(_20622__bF_buf0), .C(_19022_), .D(_20621__bF_buf0), .Y(_21616_) );
	OAI22X1 OAI22X1_645 ( .gnd(gnd), .vdd(vdd), .A(_19025_), .B(_20626__bF_buf0), .C(_19026_), .D(_20624__bF_buf0), .Y(_21617_) );
	NOR2X1 NOR2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_21617_), .B(_21616_), .Y(_21618_) );
	OAI22X1 OAI22X1_646 ( .gnd(gnd), .vdd(vdd), .A(_19029_), .B(_20629__bF_buf0), .C(_19030_), .D(_20630__bF_buf0), .Y(_21619_) );
	OAI22X1 OAI22X1_647 ( .gnd(gnd), .vdd(vdd), .A(_19033_), .B(_20633__bF_buf0), .C(_19032_), .D(_20632__bF_buf0), .Y(_21620_) );
	NOR2X1 NOR2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_21619_), .B(_21620_), .Y(_21621_) );
	NAND2X1 NAND2X1_3727 ( .gnd(gnd), .vdd(vdd), .A(_21618_), .B(_21621_), .Y(_21622_) );
	NOR2X1 NOR2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_21615_), .B(_21622_), .Y(_21623_) );
	NAND2X1 NAND2X1_3728 ( .gnd(gnd), .vdd(vdd), .A(_21623_), .B(_21609_), .Y(readB_regOut_29_) );
	NAND3X1 NAND3X1_3968 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_30_), .B(_20559__bF_buf5), .C(_20557__bF_buf2), .Y(_21624_) );
	NAND3X1 NAND3X1_3969 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_30_), .B(_20562__bF_buf5), .C(_20557__bF_buf1), .Y(_21625_) );
	NAND2X1 NAND2X1_3729 ( .gnd(gnd), .vdd(vdd), .A(_21624_), .B(_21625_), .Y(_21626_) );
	OAI22X1 OAI22X1_648 ( .gnd(gnd), .vdd(vdd), .A(_19041_), .B(_20568__bF_buf4), .C(_19042_), .D(_20567__bF_buf4), .Y(_21627_) );
	NOR2X1 NOR2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_21626_), .B(_21627_), .Y(_21628_) );
	OAI22X1 OAI22X1_649 ( .gnd(gnd), .vdd(vdd), .A(_19045_), .B(_20576__bF_buf4), .C(_19046_), .D(_20575__bF_buf4), .Y(_21629_) );
	OAI22X1 OAI22X1_650 ( .gnd(gnd), .vdd(vdd), .A(_19048_), .B(_20581__bF_buf4), .C(_19049_), .D(_20580__bF_buf4), .Y(_21630_) );
	NOR2X1 NOR2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_21630_), .B(_21629_), .Y(_21631_) );
	NAND2X1 NAND2X1_3730 ( .gnd(gnd), .vdd(vdd), .A(_21628_), .B(_21631_), .Y(_21632_) );
	OAI22X1 OAI22X1_651 ( .gnd(gnd), .vdd(vdd), .A(_19054_), .B(_20586__bF_buf4), .C(_19053_), .D(_20585__bF_buf4), .Y(_21633_) );
	NAND3X1 NAND3X1_3970 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_30_), .B(_20588__bF_buf1), .C(_20590__bF_buf3), .Y(_21634_) );
	OAI21X1 OAI21X1_4782 ( .gnd(gnd), .vdd(vdd), .A(_19056_), .B(_20589__bF_buf4), .C(_21634_), .Y(_21635_) );
	NOR2X1 NOR2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_21633_), .B(_21635_), .Y(_21636_) );
	NAND3X1 NAND3X1_3971 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_30_), .B(bLoc_frameOut_4_bF_buf6), .C(_20595__bF_buf4), .Y(_21637_) );
	OAI21X1 OAI21X1_4783 ( .gnd(gnd), .vdd(vdd), .A(_19060_), .B(_20594__bF_buf4), .C(_21637_), .Y(_21638_) );
	NAND3X1 NAND3X1_3972 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_30_), .B(_20574__bF_buf6), .C(_20590__bF_buf2), .Y(_21639_) );
	OAI21X1 OAI21X1_4784 ( .gnd(gnd), .vdd(vdd), .A(_19063_), .B(_20598__bF_buf4), .C(_21639_), .Y(_21640_) );
	NOR2X1 NOR2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_21638_), .B(_21640_), .Y(_21641_) );
	NAND2X1 NAND2X1_3731 ( .gnd(gnd), .vdd(vdd), .A(_21641_), .B(_21636_), .Y(_21642_) );
	NOR2X1 NOR2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_21642_), .B(_21632_), .Y(_21643_) );
	AOI22X1 AOI22X1_502 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf4), .B(registers_a2_30_), .C(registers_r1_30_), .D(_20606__bF_buf4), .Y(_21644_) );
	AOI22X1 AOI22X1_503 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf4), .B(registers_r4_30_), .C(registers_r5_30_), .D(_20611__bF_buf4), .Y(_21645_) );
	NAND3X1 NAND3X1_3973 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_30_), .B(_20607__bF_buf2), .C(_20574__bF_buf5), .Y(_21646_) );
	OAI21X1 OAI21X1_4785 ( .gnd(gnd), .vdd(vdd), .A(_19071_), .B(_20617__bF_buf4), .C(_21646_), .Y(_21647_) );
	AOI21X1 AOI21X1_3177 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_30_), .B(_20615__bF_buf4), .C(_21647_), .Y(_21648_) );
	NAND3X1 NAND3X1_3974 ( .gnd(gnd), .vdd(vdd), .A(_21644_), .B(_21645_), .C(_21648_), .Y(_21649_) );
	OAI22X1 OAI22X1_652 ( .gnd(gnd), .vdd(vdd), .A(_19077_), .B(_20622__bF_buf4), .C(_19076_), .D(_20621__bF_buf4), .Y(_21650_) );
	OAI22X1 OAI22X1_653 ( .gnd(gnd), .vdd(vdd), .A(_19079_), .B(_20626__bF_buf4), .C(_19080_), .D(_20624__bF_buf4), .Y(_21651_) );
	NOR2X1 NOR2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_21651_), .B(_21650_), .Y(_21652_) );
	OAI22X1 OAI22X1_654 ( .gnd(gnd), .vdd(vdd), .A(_19083_), .B(_20629__bF_buf4), .C(_19084_), .D(_20630__bF_buf4), .Y(_21653_) );
	OAI22X1 OAI22X1_655 ( .gnd(gnd), .vdd(vdd), .A(_19087_), .B(_20633__bF_buf4), .C(_19086_), .D(_20632__bF_buf4), .Y(_21654_) );
	NOR2X1 NOR2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_21653_), .B(_21654_), .Y(_21655_) );
	NAND2X1 NAND2X1_3732 ( .gnd(gnd), .vdd(vdd), .A(_21652_), .B(_21655_), .Y(_21656_) );
	NOR2X1 NOR2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_21649_), .B(_21656_), .Y(_21657_) );
	NAND2X1 NAND2X1_3733 ( .gnd(gnd), .vdd(vdd), .A(_21657_), .B(_21643_), .Y(readB_regOut_30_) );
	NAND3X1 NAND3X1_3975 ( .gnd(gnd), .vdd(vdd), .A(registers_r6_31_), .B(_20559__bF_buf4), .C(_20557__bF_buf0), .Y(_21658_) );
	NAND3X1 NAND3X1_3976 ( .gnd(gnd), .vdd(vdd), .A(registers_r7_31_), .B(_20562__bF_buf4), .C(_20557__bF_buf7), .Y(_21659_) );
	NAND2X1 NAND2X1_3734 ( .gnd(gnd), .vdd(vdd), .A(_21658_), .B(_21659_), .Y(_21660_) );
	OAI22X1 OAI22X1_656 ( .gnd(gnd), .vdd(vdd), .A(_19095_), .B(_20568__bF_buf3), .C(_19096_), .D(_20567__bF_buf3), .Y(_21661_) );
	NOR2X1 NOR2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_21660_), .B(_21661_), .Y(_21662_) );
	OAI22X1 OAI22X1_657 ( .gnd(gnd), .vdd(vdd), .A(_19099_), .B(_20576__bF_buf3), .C(_19100_), .D(_20575__bF_buf3), .Y(_21663_) );
	OAI22X1 OAI22X1_658 ( .gnd(gnd), .vdd(vdd), .A(_19102_), .B(_20581__bF_buf3), .C(_19103_), .D(_20580__bF_buf3), .Y(_21664_) );
	NOR2X1 NOR2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_21664_), .B(_21663_), .Y(_21665_) );
	NAND2X1 NAND2X1_3735 ( .gnd(gnd), .vdd(vdd), .A(_21662_), .B(_21665_), .Y(_21666_) );
	OAI22X1 OAI22X1_659 ( .gnd(gnd), .vdd(vdd), .A(_19108_), .B(_20586__bF_buf3), .C(_19107_), .D(_20585__bF_buf3), .Y(_21667_) );
	NAND3X1 NAND3X1_3977 ( .gnd(gnd), .vdd(vdd), .A(registers_r20_31_), .B(_20588__bF_buf0), .C(_20590__bF_buf1), .Y(_21668_) );
	OAI21X1 OAI21X1_4786 ( .gnd(gnd), .vdd(vdd), .A(_19110_), .B(_20589__bF_buf3), .C(_21668_), .Y(_21669_) );
	NOR2X1 NOR2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_21667_), .B(_21669_), .Y(_21670_) );
	NAND3X1 NAND3X1_3978 ( .gnd(gnd), .vdd(vdd), .A(registers_r31_31_), .B(bLoc_frameOut_4_bF_buf5), .C(_20595__bF_buf3), .Y(_21671_) );
	OAI21X1 OAI21X1_4787 ( .gnd(gnd), .vdd(vdd), .A(_19114_), .B(_20594__bF_buf3), .C(_21671_), .Y(_21672_) );
	NAND3X1 NAND3X1_3979 ( .gnd(gnd), .vdd(vdd), .A(registers_r24_31_), .B(_20574__bF_buf4), .C(_20590__bF_buf0), .Y(_21673_) );
	OAI21X1 OAI21X1_4788 ( .gnd(gnd), .vdd(vdd), .A(_19117_), .B(_20598__bF_buf3), .C(_21673_), .Y(_21674_) );
	NOR2X1 NOR2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_21672_), .B(_21674_), .Y(_21675_) );
	NAND2X1 NAND2X1_3736 ( .gnd(gnd), .vdd(vdd), .A(_21675_), .B(_21670_), .Y(_21676_) );
	NOR2X1 NOR2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_21676_), .B(_21666_), .Y(_21677_) );
	AOI22X1 AOI22X1_504 ( .gnd(gnd), .vdd(vdd), .A(_20608__bF_buf3), .B(registers_a2_31_), .C(registers_r1_31_), .D(_20606__bF_buf3), .Y(_21678_) );
	AOI22X1 AOI22X1_505 ( .gnd(gnd), .vdd(vdd), .A(_20610__bF_buf3), .B(registers_r4_31_), .C(registers_r5_31_), .D(_20611__bF_buf3), .Y(_21679_) );
	NAND3X1 NAND3X1_3980 ( .gnd(gnd), .vdd(vdd), .A(registers_fp_31_), .B(_20607__bF_buf1), .C(_20574__bF_buf3), .Y(_21680_) );
	OAI21X1 OAI21X1_4789 ( .gnd(gnd), .vdd(vdd), .A(_19125_), .B(_20617__bF_buf3), .C(_21680_), .Y(_21681_) );
	AOI21X1 AOI21X1_3178 ( .gnd(gnd), .vdd(vdd), .A(registers_a0_31_), .B(_20615__bF_buf3), .C(_21681_), .Y(_21682_) );
	NAND3X1 NAND3X1_3981 ( .gnd(gnd), .vdd(vdd), .A(_21678_), .B(_21679_), .C(_21682_), .Y(_21683_) );
	OAI22X1 OAI22X1_660 ( .gnd(gnd), .vdd(vdd), .A(_19131_), .B(_20622__bF_buf3), .C(_19130_), .D(_20621__bF_buf3), .Y(_21684_) );
	OAI22X1 OAI22X1_661 ( .gnd(gnd), .vdd(vdd), .A(_19133_), .B(_20626__bF_buf3), .C(_19134_), .D(_20624__bF_buf3), .Y(_21685_) );
	NOR2X1 NOR2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_21685_), .B(_21684_), .Y(_21686_) );
	OAI22X1 OAI22X1_662 ( .gnd(gnd), .vdd(vdd), .A(_19137_), .B(_20629__bF_buf3), .C(_19138_), .D(_20630__bF_buf3), .Y(_21687_) );
	OAI22X1 OAI22X1_663 ( .gnd(gnd), .vdd(vdd), .A(_19141_), .B(_20633__bF_buf3), .C(_19140_), .D(_20632__bF_buf3), .Y(_21688_) );
	NOR2X1 NOR2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_21687_), .B(_21688_), .Y(_21689_) );
	NAND2X1 NAND2X1_3737 ( .gnd(gnd), .vdd(vdd), .A(_21686_), .B(_21689_), .Y(_21690_) );
	NOR2X1 NOR2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_21683_), .B(_21690_), .Y(_21691_) );
	NAND2X1 NAND2X1_3738 ( .gnd(gnd), .vdd(vdd), .A(_21691_), .B(_21677_), .Y(readB_regOut_31_) );
	DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17349__0_), .Q(registers_r1_0_) );
	DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17349__1_), .Q(registers_r1_1_) );
	DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17349__2_), .Q(registers_r1_2_) );
	DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17349__3_), .Q(registers_r1_3_) );
	DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17349__4_), .Q(registers_r1_4_) );
	DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17349__5_), .Q(registers_r1_5_) );
	DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17349__6_), .Q(registers_r1_6_) );
	DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17349__7_), .Q(registers_r1_7_) );
	DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17349__8_), .Q(registers_r1_8_) );
	DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17349__9_), .Q(registers_r1_9_) );
	DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17349__10_), .Q(registers_r1_10_) );
	DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17349__11_), .Q(registers_r1_11_) );
	DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17349__12_), .Q(registers_r1_12_) );
	DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17349__13_), .Q(registers_r1_13_) );
	DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17349__14_), .Q(registers_r1_14_) );
	DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17349__15_), .Q(registers_r1_15_) );
	DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17349__16_), .Q(registers_r1_16_) );
	DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17349__17_), .Q(registers_r1_17_) );
	DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17349__18_), .Q(registers_r1_18_) );
	DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17349__19_), .Q(registers_r1_19_) );
	DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17349__20_), .Q(registers_r1_20_) );
	DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17349__21_), .Q(registers_r1_21_) );
	DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17349__22_), .Q(registers_r1_22_) );
	DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17349__23_), .Q(registers_r1_23_) );
	DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17349__24_), .Q(registers_r1_24_) );
	DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17349__25_), .Q(registers_r1_25_) );
	DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17349__26_), .Q(registers_r1_26_) );
	DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17349__27_), .Q(registers_r1_27_) );
	DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17349__28_), .Q(registers_r1_28_) );
	DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17349__29_), .Q(registers_r1_29_) );
	DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17349__30_), .Q(registers_r1_30_) );
	DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17349__31_), .Q(registers_r1_31_) );
	DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17360__0_), .Q(registers_r2_0_) );
	DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17360__1_), .Q(registers_r2_1_) );
	DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17360__2_), .Q(registers_r2_2_) );
	DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17360__3_), .Q(registers_r2_3_) );
	DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17360__4_), .Q(registers_r2_4_) );
	DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17360__5_), .Q(registers_r2_5_) );
	DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17360__6_), .Q(registers_r2_6_) );
	DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17360__7_), .Q(registers_r2_7_) );
	DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17360__8_), .Q(registers_r2_8_) );
	DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17360__9_), .Q(registers_r2_9_) );
	DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17360__10_), .Q(registers_r2_10_) );
	DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17360__11_), .Q(registers_r2_11_) );
	DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17360__12_), .Q(registers_r2_12_) );
	DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17360__13_), .Q(registers_r2_13_) );
	DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17360__14_), .Q(registers_r2_14_) );
	DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17360__15_), .Q(registers_r2_15_) );
	DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17360__16_), .Q(registers_r2_16_) );
	DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17360__17_), .Q(registers_r2_17_) );
	DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17360__18_), .Q(registers_r2_18_) );
	DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17360__19_), .Q(registers_r2_19_) );
	DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17360__20_), .Q(registers_r2_20_) );
	DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17360__21_), .Q(registers_r2_21_) );
	DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17360__22_), .Q(registers_r2_22_) );
	DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17360__23_), .Q(registers_r2_23_) );
	DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17360__24_), .Q(registers_r2_24_) );
	DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17360__25_), .Q(registers_r2_25_) );
	DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17360__26_), .Q(registers_r2_26_) );
	DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17360__27_), .Q(registers_r2_27_) );
	DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17360__28_), .Q(registers_r2_28_) );
	DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17360__29_), .Q(registers_r2_29_) );
	DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17360__30_), .Q(registers_r2_30_) );
	DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17360__31_), .Q(registers_r2_31_) );
	DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17363__0_), .Q(registers_gp_0_) );
	DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17363__1_), .Q(registers_gp_1_) );
	DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17363__2_), .Q(registers_gp_2_) );
	DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17363__3_), .Q(registers_gp_3_) );
	DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17363__4_), .Q(registers_gp_4_) );
	DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17363__5_), .Q(registers_gp_5_) );
	DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17363__6_), .Q(registers_gp_6_) );
	DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17363__7_), .Q(registers_gp_7_) );
	DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17363__8_), .Q(registers_gp_8_) );
	DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17363__9_), .Q(registers_gp_9_) );
	DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17363__10_), .Q(registers_gp_10_) );
	DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17363__11_), .Q(registers_gp_11_) );
	DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17363__12_), .Q(registers_gp_12_) );
	DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17363__13_), .Q(registers_gp_13_) );
	DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17363__14_), .Q(registers_gp_14_) );
	DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17363__15_), .Q(registers_gp_15_) );
	DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17363__16_), .Q(registers_gp_16_) );
	DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17363__17_), .Q(registers_gp_17_) );
	DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17363__18_), .Q(registers_gp_18_) );
	DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17363__19_), .Q(registers_gp_19_) );
	DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17363__20_), .Q(registers_gp_20_) );
	DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17363__21_), .Q(registers_gp_21_) );
	DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17363__22_), .Q(registers_gp_22_) );
	DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17363__23_), .Q(registers_gp_23_) );
	DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17363__24_), .Q(registers_gp_24_) );
	DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17363__25_), .Q(registers_gp_25_) );
	DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17363__26_), .Q(registers_gp_26_) );
	DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17363__27_), .Q(registers_gp_27_) );
	DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17363__28_), .Q(registers_gp_28_) );
	DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17363__29_), .Q(registers_gp_29_) );
	DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17363__30_), .Q(registers_gp_30_) );
	DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17363__31_), .Q(registers_gp_31_) );
	DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17364__0_), .Q(registers_r4_0_) );
	DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17364__1_), .Q(registers_r4_1_) );
	DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17364__2_), .Q(registers_r4_2_) );
	DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17364__3_), .Q(registers_r4_3_) );
	DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17364__4_), .Q(registers_r4_4_) );
	DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17364__5_), .Q(registers_r4_5_) );
	DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17364__6_), .Q(registers_r4_6_) );
	DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17364__7_), .Q(registers_r4_7_) );
	DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17364__8_), .Q(registers_r4_8_) );
	DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17364__9_), .Q(registers_r4_9_) );
	DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17364__10_), .Q(registers_r4_10_) );
	DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17364__11_), .Q(registers_r4_11_) );
	DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17364__12_), .Q(registers_r4_12_) );
	DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17364__13_), .Q(registers_r4_13_) );
	DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17364__14_), .Q(registers_r4_14_) );
	DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17364__15_), .Q(registers_r4_15_) );
	DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17364__16_), .Q(registers_r4_16_) );
	DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17364__17_), .Q(registers_r4_17_) );
	DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17364__18_), .Q(registers_r4_18_) );
	DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17364__19_), .Q(registers_r4_19_) );
	DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17364__20_), .Q(registers_r4_20_) );
	DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17364__21_), .Q(registers_r4_21_) );
	DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17364__22_), .Q(registers_r4_22_) );
	DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17364__23_), .Q(registers_r4_23_) );
	DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17364__24_), .Q(registers_r4_24_) );
	DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17364__25_), .Q(registers_r4_25_) );
	DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17364__26_), .Q(registers_r4_26_) );
	DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17364__27_), .Q(registers_r4_27_) );
	DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17364__28_), .Q(registers_r4_28_) );
	DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17364__29_), .Q(registers_r4_29_) );
	DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17364__30_), .Q(registers_r4_30_) );
	DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17364__31_), .Q(registers_r4_31_) );
	DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17365__0_), .Q(registers_r5_0_) );
	DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17365__1_), .Q(registers_r5_1_) );
	DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17365__2_), .Q(registers_r5_2_) );
	DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17365__3_), .Q(registers_r5_3_) );
	DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17365__4_), .Q(registers_r5_4_) );
	DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17365__5_), .Q(registers_r5_5_) );
	DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17365__6_), .Q(registers_r5_6_) );
	DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17365__7_), .Q(registers_r5_7_) );
	DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17365__8_), .Q(registers_r5_8_) );
	DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17365__9_), .Q(registers_r5_9_) );
	DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17365__10_), .Q(registers_r5_10_) );
	DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17365__11_), .Q(registers_r5_11_) );
	DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17365__12_), .Q(registers_r5_12_) );
	DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17365__13_), .Q(registers_r5_13_) );
	DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17365__14_), .Q(registers_r5_14_) );
	DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17365__15_), .Q(registers_r5_15_) );
	DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17365__16_), .Q(registers_r5_16_) );
	DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17365__17_), .Q(registers_r5_17_) );
	DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17365__18_), .Q(registers_r5_18_) );
	DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17365__19_), .Q(registers_r5_19_) );
	DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17365__20_), .Q(registers_r5_20_) );
	DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17365__21_), .Q(registers_r5_21_) );
	DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17365__22_), .Q(registers_r5_22_) );
	DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17365__23_), .Q(registers_r5_23_) );
	DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17365__24_), .Q(registers_r5_24_) );
	DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17365__25_), .Q(registers_r5_25_) );
	DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17365__26_), .Q(registers_r5_26_) );
	DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17365__27_), .Q(registers_r5_27_) );
	DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17365__28_), .Q(registers_r5_28_) );
	DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17365__29_), .Q(registers_r5_29_) );
	DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17365__30_), .Q(registers_r5_30_) );
	DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17365__31_), .Q(registers_r5_31_) );
	DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17366__0_), .Q(registers_r6_0_) );
	DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17366__1_), .Q(registers_r6_1_) );
	DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17366__2_), .Q(registers_r6_2_) );
	DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17366__3_), .Q(registers_r6_3_) );
	DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17366__4_), .Q(registers_r6_4_) );
	DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17366__5_), .Q(registers_r6_5_) );
	DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17366__6_), .Q(registers_r6_6_) );
	DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17366__7_), .Q(registers_r6_7_) );
	DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17366__8_), .Q(registers_r6_8_) );
	DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17366__9_), .Q(registers_r6_9_) );
	DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17366__10_), .Q(registers_r6_10_) );
	DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17366__11_), .Q(registers_r6_11_) );
	DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17366__12_), .Q(registers_r6_12_) );
	DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17366__13_), .Q(registers_r6_13_) );
	DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17366__14_), .Q(registers_r6_14_) );
	DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17366__15_), .Q(registers_r6_15_) );
	DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17366__16_), .Q(registers_r6_16_) );
	DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17366__17_), .Q(registers_r6_17_) );
	DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17366__18_), .Q(registers_r6_18_) );
	DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17366__19_), .Q(registers_r6_19_) );
	DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17366__20_), .Q(registers_r6_20_) );
	DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17366__21_), .Q(registers_r6_21_) );
	DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17366__22_), .Q(registers_r6_22_) );
	DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17366__23_), .Q(registers_r6_23_) );
	DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17366__24_), .Q(registers_r6_24_) );
	DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17366__25_), .Q(registers_r6_25_) );
	DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17366__26_), .Q(registers_r6_26_) );
	DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17366__27_), .Q(registers_r6_27_) );
	DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17366__28_), .Q(registers_r6_28_) );
	DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17366__29_), .Q(registers_r6_29_) );
	DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17366__30_), .Q(registers_r6_30_) );
	DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17366__31_), .Q(registers_r6_31_) );
	DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17367__0_), .Q(registers_r7_0_) );
	DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17367__1_), .Q(registers_r7_1_) );
	DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17367__2_), .Q(registers_r7_2_) );
	DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17367__3_), .Q(registers_r7_3_) );
	DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17367__4_), .Q(registers_r7_4_) );
	DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17367__5_), .Q(registers_r7_5_) );
	DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17367__6_), .Q(registers_r7_6_) );
	DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17367__7_), .Q(registers_r7_7_) );
	DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17367__8_), .Q(registers_r7_8_) );
	DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17367__9_), .Q(registers_r7_9_) );
	DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17367__10_), .Q(registers_r7_10_) );
	DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17367__11_), .Q(registers_r7_11_) );
	DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17367__12_), .Q(registers_r7_12_) );
	DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17367__13_), .Q(registers_r7_13_) );
	DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17367__14_), .Q(registers_r7_14_) );
	DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17367__15_), .Q(registers_r7_15_) );
	DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17367__16_), .Q(registers_r7_16_) );
	DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17367__17_), .Q(registers_r7_17_) );
	DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17367__18_), .Q(registers_r7_18_) );
	DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17367__19_), .Q(registers_r7_19_) );
	DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17367__20_), .Q(registers_r7_20_) );
	DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17367__21_), .Q(registers_r7_21_) );
	DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17367__22_), .Q(registers_r7_22_) );
	DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17367__23_), .Q(registers_r7_23_) );
	DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17367__24_), .Q(registers_r7_24_) );
	DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17367__25_), .Q(registers_r7_25_) );
	DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17367__26_), .Q(registers_r7_26_) );
	DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17367__27_), .Q(registers_r7_27_) );
	DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17367__28_), .Q(registers_r7_28_) );
	DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17367__29_), .Q(registers_r7_29_) );
	DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17367__30_), .Q(registers_r7_30_) );
	DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17367__31_), .Q(registers_r7_31_) );
	DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17368__0_), .Q(registers_fp_0_) );
	DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17368__1_), .Q(registers_fp_1_) );
	DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17368__2_), .Q(registers_fp_2_) );
	DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17368__3_), .Q(registers_fp_3_) );
	DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17368__4_), .Q(registers_fp_4_) );
	DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17368__5_), .Q(registers_fp_5_) );
	DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17368__6_), .Q(registers_fp_6_) );
	DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17368__7_), .Q(registers_fp_7_) );
	DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17368__8_), .Q(registers_fp_8_) );
	DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17368__9_), .Q(registers_fp_9_) );
	DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17368__10_), .Q(registers_fp_10_) );
	DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17368__11_), .Q(registers_fp_11_) );
	DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17368__12_), .Q(registers_fp_12_) );
	DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17368__13_), .Q(registers_fp_13_) );
	DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17368__14_), .Q(registers_fp_14_) );
	DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17368__15_), .Q(registers_fp_15_) );
	DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17368__16_), .Q(registers_fp_16_) );
	DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17368__17_), .Q(registers_fp_17_) );
	DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17368__18_), .Q(registers_fp_18_) );
	DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17368__19_), .Q(registers_fp_19_) );
	DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17368__20_), .Q(registers_fp_20_) );
	DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17368__21_), .Q(registers_fp_21_) );
	DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17368__22_), .Q(registers_fp_22_) );
	DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17368__23_), .Q(registers_fp_23_) );
	DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17368__24_), .Q(registers_fp_24_) );
	DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17368__25_), .Q(registers_fp_25_) );
	DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17368__26_), .Q(registers_fp_26_) );
	DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17368__27_), .Q(registers_fp_27_) );
	DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17368__28_), .Q(registers_fp_28_) );
	DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17368__29_), .Q(registers_fp_29_) );
	DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17368__30_), .Q(registers_fp_30_) );
	DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17368__31_), .Q(registers_fp_31_) );
	DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17369__0_), .Q(registers_r9_0_) );
	DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17369__1_), .Q(registers_r9_1_) );
	DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17369__2_), .Q(registers_r9_2_) );
	DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17369__3_), .Q(registers_r9_3_) );
	DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17369__4_), .Q(registers_r9_4_) );
	DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17369__5_), .Q(registers_r9_5_) );
	DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17369__6_), .Q(registers_r9_6_) );
	DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17369__7_), .Q(registers_r9_7_) );
	DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17369__8_), .Q(registers_r9_8_) );
	DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17369__9_), .Q(registers_r9_9_) );
	DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17369__10_), .Q(registers_r9_10_) );
	DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17369__11_), .Q(registers_r9_11_) );
	DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17369__12_), .Q(registers_r9_12_) );
	DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17369__13_), .Q(registers_r9_13_) );
	DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17369__14_), .Q(registers_r9_14_) );
	DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17369__15_), .Q(registers_r9_15_) );
	DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17369__16_), .Q(registers_r9_16_) );
	DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17369__17_), .Q(registers_r9_17_) );
	DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17369__18_), .Q(registers_r9_18_) );
	DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17369__19_), .Q(registers_r9_19_) );
	DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17369__20_), .Q(registers_r9_20_) );
	DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17369__21_), .Q(registers_r9_21_) );
	DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17369__22_), .Q(registers_r9_22_) );
	DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17369__23_), .Q(registers_r9_23_) );
	DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17369__24_), .Q(registers_r9_24_) );
	DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17369__25_), .Q(registers_r9_25_) );
	DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17369__26_), .Q(registers_r9_26_) );
	DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17369__27_), .Q(registers_r9_27_) );
	DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17369__28_), .Q(registers_r9_28_) );
	DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17369__29_), .Q(registers_r9_29_) );
	DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17369__30_), .Q(registers_r9_30_) );
	DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17369__31_), .Q(registers_r9_31_) );
	DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17339__0_), .Q(registers_a0_0_) );
	DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17339__1_), .Q(registers_a0_1_) );
	DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17339__2_), .Q(registers_a0_2_) );
	DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17339__3_), .Q(registers_a0_3_) );
	DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17339__4_), .Q(registers_a0_4_) );
	DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17339__5_), .Q(registers_a0_5_) );
	DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17339__6_), .Q(registers_a0_6_) );
	DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17339__7_), .Q(registers_a0_7_) );
	DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17339__8_), .Q(registers_a0_8_) );
	DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17339__9_), .Q(registers_a0_9_) );
	DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17339__10_), .Q(registers_a0_10_) );
	DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17339__11_), .Q(registers_a0_11_) );
	DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17339__12_), .Q(registers_a0_12_) );
	DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17339__13_), .Q(registers_a0_13_) );
	DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17339__14_), .Q(registers_a0_14_) );
	DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17339__15_), .Q(registers_a0_15_) );
	DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17339__16_), .Q(registers_a0_16_) );
	DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17339__17_), .Q(registers_a0_17_) );
	DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17339__18_), .Q(registers_a0_18_) );
	DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17339__19_), .Q(registers_a0_19_) );
	DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17339__20_), .Q(registers_a0_20_) );
	DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17339__21_), .Q(registers_a0_21_) );
	DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17339__22_), .Q(registers_a0_22_) );
	DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17339__23_), .Q(registers_a0_23_) );
	DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17339__24_), .Q(registers_a0_24_) );
	DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17339__25_), .Q(registers_a0_25_) );
	DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17339__26_), .Q(registers_a0_26_) );
	DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17339__27_), .Q(registers_a0_27_) );
	DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17339__28_), .Q(registers_a0_28_) );
	DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17339__29_), .Q(registers_a0_29_) );
	DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17339__30_), .Q(registers_a0_30_) );
	DFFPOSX1 DFFPOSX1_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17339__31_), .Q(registers_a0_31_) );
	DFFPOSX1 DFFPOSX1_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17340__0_), .Q(registers_a1_0_) );
	DFFPOSX1 DFFPOSX1_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17340__1_), .Q(registers_a1_1_) );
	DFFPOSX1 DFFPOSX1_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17340__2_), .Q(registers_a1_2_) );
	DFFPOSX1 DFFPOSX1_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17340__3_), .Q(registers_a1_3_) );
	DFFPOSX1 DFFPOSX1_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17340__4_), .Q(registers_a1_4_) );
	DFFPOSX1 DFFPOSX1_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17340__5_), .Q(registers_a1_5_) );
	DFFPOSX1 DFFPOSX1_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17340__6_), .Q(registers_a1_6_) );
	DFFPOSX1 DFFPOSX1_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17340__7_), .Q(registers_a1_7_) );
	DFFPOSX1 DFFPOSX1_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17340__8_), .Q(registers_a1_8_) );
	DFFPOSX1 DFFPOSX1_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17340__9_), .Q(registers_a1_9_) );
	DFFPOSX1 DFFPOSX1_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17340__10_), .Q(registers_a1_10_) );
	DFFPOSX1 DFFPOSX1_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17340__11_), .Q(registers_a1_11_) );
	DFFPOSX1 DFFPOSX1_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17340__12_), .Q(registers_a1_12_) );
	DFFPOSX1 DFFPOSX1_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17340__13_), .Q(registers_a1_13_) );
	DFFPOSX1 DFFPOSX1_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17340__14_), .Q(registers_a1_14_) );
	DFFPOSX1 DFFPOSX1_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17340__15_), .Q(registers_a1_15_) );
	DFFPOSX1 DFFPOSX1_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17340__16_), .Q(registers_a1_16_) );
	DFFPOSX1 DFFPOSX1_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17340__17_), .Q(registers_a1_17_) );
	DFFPOSX1 DFFPOSX1_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17340__18_), .Q(registers_a1_18_) );
	DFFPOSX1 DFFPOSX1_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17340__19_), .Q(registers_a1_19_) );
	DFFPOSX1 DFFPOSX1_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17340__20_), .Q(registers_a1_20_) );
	DFFPOSX1 DFFPOSX1_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17340__21_), .Q(registers_a1_21_) );
	DFFPOSX1 DFFPOSX1_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17340__22_), .Q(registers_a1_22_) );
	DFFPOSX1 DFFPOSX1_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17340__23_), .Q(registers_a1_23_) );
	DFFPOSX1 DFFPOSX1_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17340__24_), .Q(registers_a1_24_) );
	DFFPOSX1 DFFPOSX1_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17340__25_), .Q(registers_a1_25_) );
	DFFPOSX1 DFFPOSX1_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17340__26_), .Q(registers_a1_26_) );
	DFFPOSX1 DFFPOSX1_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17340__27_), .Q(registers_a1_27_) );
	DFFPOSX1 DFFPOSX1_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17340__28_), .Q(registers_a1_28_) );
	DFFPOSX1 DFFPOSX1_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17340__29_), .Q(registers_a1_29_) );
	DFFPOSX1 DFFPOSX1_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17340__30_), .Q(registers_a1_30_) );
	DFFPOSX1 DFFPOSX1_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17340__31_), .Q(registers_a1_31_) );
	DFFPOSX1 DFFPOSX1_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17341__0_), .Q(registers_a2_0_) );
	DFFPOSX1 DFFPOSX1_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17341__1_), .Q(registers_a2_1_) );
	DFFPOSX1 DFFPOSX1_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17341__2_), .Q(registers_a2_2_) );
	DFFPOSX1 DFFPOSX1_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17341__3_), .Q(registers_a2_3_) );
	DFFPOSX1 DFFPOSX1_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17341__4_), .Q(registers_a2_4_) );
	DFFPOSX1 DFFPOSX1_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17341__5_), .Q(registers_a2_5_) );
	DFFPOSX1 DFFPOSX1_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17341__6_), .Q(registers_a2_6_) );
	DFFPOSX1 DFFPOSX1_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17341__7_), .Q(registers_a2_7_) );
	DFFPOSX1 DFFPOSX1_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17341__8_), .Q(registers_a2_8_) );
	DFFPOSX1 DFFPOSX1_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17341__9_), .Q(registers_a2_9_) );
	DFFPOSX1 DFFPOSX1_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17341__10_), .Q(registers_a2_10_) );
	DFFPOSX1 DFFPOSX1_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17341__11_), .Q(registers_a2_11_) );
	DFFPOSX1 DFFPOSX1_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17341__12_), .Q(registers_a2_12_) );
	DFFPOSX1 DFFPOSX1_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17341__13_), .Q(registers_a2_13_) );
	DFFPOSX1 DFFPOSX1_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17341__14_), .Q(registers_a2_14_) );
	DFFPOSX1 DFFPOSX1_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17341__15_), .Q(registers_a2_15_) );
	DFFPOSX1 DFFPOSX1_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17341__16_), .Q(registers_a2_16_) );
	DFFPOSX1 DFFPOSX1_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17341__17_), .Q(registers_a2_17_) );
	DFFPOSX1 DFFPOSX1_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17341__18_), .Q(registers_a2_18_) );
	DFFPOSX1 DFFPOSX1_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17341__19_), .Q(registers_a2_19_) );
	DFFPOSX1 DFFPOSX1_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17341__20_), .Q(registers_a2_20_) );
	DFFPOSX1 DFFPOSX1_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17341__21_), .Q(registers_a2_21_) );
	DFFPOSX1 DFFPOSX1_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17341__22_), .Q(registers_a2_22_) );
	DFFPOSX1 DFFPOSX1_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17341__23_), .Q(registers_a2_23_) );
	DFFPOSX1 DFFPOSX1_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17341__24_), .Q(registers_a2_24_) );
	DFFPOSX1 DFFPOSX1_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17341__25_), .Q(registers_a2_25_) );
	DFFPOSX1 DFFPOSX1_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17341__26_), .Q(registers_a2_26_) );
	DFFPOSX1 DFFPOSX1_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17341__27_), .Q(registers_a2_27_) );
	DFFPOSX1 DFFPOSX1_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17341__28_), .Q(registers_a2_28_) );
	DFFPOSX1 DFFPOSX1_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17341__29_), .Q(registers_a2_29_) );
	DFFPOSX1 DFFPOSX1_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17341__30_), .Q(registers_a2_30_) );
	DFFPOSX1 DFFPOSX1_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17341__31_), .Q(registers_a2_31_) );
	DFFPOSX1 DFFPOSX1_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17342__0_), .Q(registers_a3_0_) );
	DFFPOSX1 DFFPOSX1_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17342__1_), .Q(registers_a3_1_) );
	DFFPOSX1 DFFPOSX1_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17342__2_), .Q(registers_a3_2_) );
	DFFPOSX1 DFFPOSX1_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17342__3_), .Q(registers_a3_3_) );
	DFFPOSX1 DFFPOSX1_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17342__4_), .Q(registers_a3_4_) );
	DFFPOSX1 DFFPOSX1_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17342__5_), .Q(registers_a3_5_) );
	DFFPOSX1 DFFPOSX1_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17342__6_), .Q(registers_a3_6_) );
	DFFPOSX1 DFFPOSX1_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17342__7_), .Q(registers_a3_7_) );
	DFFPOSX1 DFFPOSX1_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17342__8_), .Q(registers_a3_8_) );
	DFFPOSX1 DFFPOSX1_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17342__9_), .Q(registers_a3_9_) );
	DFFPOSX1 DFFPOSX1_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17342__10_), .Q(registers_a3_10_) );
	DFFPOSX1 DFFPOSX1_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17342__11_), .Q(registers_a3_11_) );
	DFFPOSX1 DFFPOSX1_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17342__12_), .Q(registers_a3_12_) );
	DFFPOSX1 DFFPOSX1_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17342__13_), .Q(registers_a3_13_) );
	DFFPOSX1 DFFPOSX1_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17342__14_), .Q(registers_a3_14_) );
	DFFPOSX1 DFFPOSX1_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17342__15_), .Q(registers_a3_15_) );
	DFFPOSX1 DFFPOSX1_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17342__16_), .Q(registers_a3_16_) );
	DFFPOSX1 DFFPOSX1_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17342__17_), .Q(registers_a3_17_) );
	DFFPOSX1 DFFPOSX1_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17342__18_), .Q(registers_a3_18_) );
	DFFPOSX1 DFFPOSX1_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17342__19_), .Q(registers_a3_19_) );
	DFFPOSX1 DFFPOSX1_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17342__20_), .Q(registers_a3_20_) );
	DFFPOSX1 DFFPOSX1_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17342__21_), .Q(registers_a3_21_) );
	DFFPOSX1 DFFPOSX1_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17342__22_), .Q(registers_a3_22_) );
	DFFPOSX1 DFFPOSX1_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17342__23_), .Q(registers_a3_23_) );
	DFFPOSX1 DFFPOSX1_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17342__24_), .Q(registers_a3_24_) );
	DFFPOSX1 DFFPOSX1_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17342__25_), .Q(registers_a3_25_) );
	DFFPOSX1 DFFPOSX1_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17342__26_), .Q(registers_a3_26_) );
	DFFPOSX1 DFFPOSX1_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17342__27_), .Q(registers_a3_27_) );
	DFFPOSX1 DFFPOSX1_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17342__28_), .Q(registers_a3_28_) );
	DFFPOSX1 DFFPOSX1_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17342__29_), .Q(registers_a3_29_) );
	DFFPOSX1 DFFPOSX1_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17342__30_), .Q(registers_a3_30_) );
	DFFPOSX1 DFFPOSX1_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17342__31_), .Q(registers_a3_31_) );
	DFFPOSX1 DFFPOSX1_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17343__0_), .Q(registers_a4_0_) );
	DFFPOSX1 DFFPOSX1_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17343__1_), .Q(registers_a4_1_) );
	DFFPOSX1 DFFPOSX1_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17343__2_), .Q(registers_a4_2_) );
	DFFPOSX1 DFFPOSX1_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17343__3_), .Q(registers_a4_3_) );
	DFFPOSX1 DFFPOSX1_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17343__4_), .Q(registers_a4_4_) );
	DFFPOSX1 DFFPOSX1_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17343__5_), .Q(registers_a4_5_) );
	DFFPOSX1 DFFPOSX1_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17343__6_), .Q(registers_a4_6_) );
	DFFPOSX1 DFFPOSX1_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17343__7_), .Q(registers_a4_7_) );
	DFFPOSX1 DFFPOSX1_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17343__8_), .Q(registers_a4_8_) );
	DFFPOSX1 DFFPOSX1_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17343__9_), .Q(registers_a4_9_) );
	DFFPOSX1 DFFPOSX1_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17343__10_), .Q(registers_a4_10_) );
	DFFPOSX1 DFFPOSX1_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17343__11_), .Q(registers_a4_11_) );
	DFFPOSX1 DFFPOSX1_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17343__12_), .Q(registers_a4_12_) );
	DFFPOSX1 DFFPOSX1_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17343__13_), .Q(registers_a4_13_) );
	DFFPOSX1 DFFPOSX1_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17343__14_), .Q(registers_a4_14_) );
	DFFPOSX1 DFFPOSX1_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17343__15_), .Q(registers_a4_15_) );
	DFFPOSX1 DFFPOSX1_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17343__16_), .Q(registers_a4_16_) );
	DFFPOSX1 DFFPOSX1_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17343__17_), .Q(registers_a4_17_) );
	DFFPOSX1 DFFPOSX1_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17343__18_), .Q(registers_a4_18_) );
	DFFPOSX1 DFFPOSX1_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17343__19_), .Q(registers_a4_19_) );
	DFFPOSX1 DFFPOSX1_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17343__20_), .Q(registers_a4_20_) );
	DFFPOSX1 DFFPOSX1_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17343__21_), .Q(registers_a4_21_) );
	DFFPOSX1 DFFPOSX1_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17343__22_), .Q(registers_a4_22_) );
	DFFPOSX1 DFFPOSX1_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17343__23_), .Q(registers_a4_23_) );
	DFFPOSX1 DFFPOSX1_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17343__24_), .Q(registers_a4_24_) );
	DFFPOSX1 DFFPOSX1_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17343__25_), .Q(registers_a4_25_) );
	DFFPOSX1 DFFPOSX1_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17343__26_), .Q(registers_a4_26_) );
	DFFPOSX1 DFFPOSX1_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17343__27_), .Q(registers_a4_27_) );
	DFFPOSX1 DFFPOSX1_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17343__28_), .Q(registers_a4_28_) );
	DFFPOSX1 DFFPOSX1_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17343__29_), .Q(registers_a4_29_) );
	DFFPOSX1 DFFPOSX1_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17343__30_), .Q(registers_a4_30_) );
	DFFPOSX1 DFFPOSX1_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17343__31_), .Q(registers_a4_31_) );
	DFFPOSX1 DFFPOSX1_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17344__0_), .Q(registers_a5_0_) );
	DFFPOSX1 DFFPOSX1_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17344__1_), .Q(registers_a5_1_) );
	DFFPOSX1 DFFPOSX1_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17344__2_), .Q(registers_a5_2_) );
	DFFPOSX1 DFFPOSX1_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17344__3_), .Q(registers_a5_3_) );
	DFFPOSX1 DFFPOSX1_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17344__4_), .Q(registers_a5_4_) );
	DFFPOSX1 DFFPOSX1_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17344__5_), .Q(registers_a5_5_) );
	DFFPOSX1 DFFPOSX1_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17344__6_), .Q(registers_a5_6_) );
	DFFPOSX1 DFFPOSX1_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17344__7_), .Q(registers_a5_7_) );
	DFFPOSX1 DFFPOSX1_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17344__8_), .Q(registers_a5_8_) );
	DFFPOSX1 DFFPOSX1_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17344__9_), .Q(registers_a5_9_) );
	DFFPOSX1 DFFPOSX1_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17344__10_), .Q(registers_a5_10_) );
	DFFPOSX1 DFFPOSX1_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17344__11_), .Q(registers_a5_11_) );
	DFFPOSX1 DFFPOSX1_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17344__12_), .Q(registers_a5_12_) );
	DFFPOSX1 DFFPOSX1_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17344__13_), .Q(registers_a5_13_) );
	DFFPOSX1 DFFPOSX1_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17344__14_), .Q(registers_a5_14_) );
	DFFPOSX1 DFFPOSX1_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17344__15_), .Q(registers_a5_15_) );
	DFFPOSX1 DFFPOSX1_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17344__16_), .Q(registers_a5_16_) );
	DFFPOSX1 DFFPOSX1_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17344__17_), .Q(registers_a5_17_) );
	DFFPOSX1 DFFPOSX1_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17344__18_), .Q(registers_a5_18_) );
	DFFPOSX1 DFFPOSX1_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17344__19_), .Q(registers_a5_19_) );
	DFFPOSX1 DFFPOSX1_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17344__20_), .Q(registers_a5_20_) );
	DFFPOSX1 DFFPOSX1_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17344__21_), .Q(registers_a5_21_) );
	DFFPOSX1 DFFPOSX1_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17344__22_), .Q(registers_a5_22_) );
	DFFPOSX1 DFFPOSX1_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17344__23_), .Q(registers_a5_23_) );
	DFFPOSX1 DFFPOSX1_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17344__24_), .Q(registers_a5_24_) );
	DFFPOSX1 DFFPOSX1_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17344__25_), .Q(registers_a5_25_) );
	DFFPOSX1 DFFPOSX1_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17344__26_), .Q(registers_a5_26_) );
	DFFPOSX1 DFFPOSX1_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17344__27_), .Q(registers_a5_27_) );
	DFFPOSX1 DFFPOSX1_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17344__28_), .Q(registers_a5_28_) );
	DFFPOSX1 DFFPOSX1_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17344__29_), .Q(registers_a5_29_) );
	DFFPOSX1 DFFPOSX1_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17344__30_), .Q(registers_a5_30_) );
	DFFPOSX1 DFFPOSX1_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17344__31_), .Q(registers_a5_31_) );
	DFFPOSX1 DFFPOSX1_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17345__0_), .Q(registers_a6_0_) );
	DFFPOSX1 DFFPOSX1_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17345__1_), .Q(registers_a6_1_) );
	DFFPOSX1 DFFPOSX1_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17345__2_), .Q(registers_a6_2_) );
	DFFPOSX1 DFFPOSX1_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17345__3_), .Q(registers_a6_3_) );
	DFFPOSX1 DFFPOSX1_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17345__4_), .Q(registers_a6_4_) );
	DFFPOSX1 DFFPOSX1_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17345__5_), .Q(registers_a6_5_) );
	DFFPOSX1 DFFPOSX1_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17345__6_), .Q(registers_a6_6_) );
	DFFPOSX1 DFFPOSX1_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17345__7_), .Q(registers_a6_7_) );
	DFFPOSX1 DFFPOSX1_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17345__8_), .Q(registers_a6_8_) );
	DFFPOSX1 DFFPOSX1_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17345__9_), .Q(registers_a6_9_) );
	DFFPOSX1 DFFPOSX1_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17345__10_), .Q(registers_a6_10_) );
	DFFPOSX1 DFFPOSX1_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17345__11_), .Q(registers_a6_11_) );
	DFFPOSX1 DFFPOSX1_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17345__12_), .Q(registers_a6_12_) );
	DFFPOSX1 DFFPOSX1_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17345__13_), .Q(registers_a6_13_) );
	DFFPOSX1 DFFPOSX1_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17345__14_), .Q(registers_a6_14_) );
	DFFPOSX1 DFFPOSX1_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17345__15_), .Q(registers_a6_15_) );
	DFFPOSX1 DFFPOSX1_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17345__16_), .Q(registers_a6_16_) );
	DFFPOSX1 DFFPOSX1_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17345__17_), .Q(registers_a6_17_) );
	DFFPOSX1 DFFPOSX1_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17345__18_), .Q(registers_a6_18_) );
	DFFPOSX1 DFFPOSX1_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17345__19_), .Q(registers_a6_19_) );
	DFFPOSX1 DFFPOSX1_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17345__20_), .Q(registers_a6_20_) );
	DFFPOSX1 DFFPOSX1_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17345__21_), .Q(registers_a6_21_) );
	DFFPOSX1 DFFPOSX1_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17345__22_), .Q(registers_a6_22_) );
	DFFPOSX1 DFFPOSX1_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17345__23_), .Q(registers_a6_23_) );
	DFFPOSX1 DFFPOSX1_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17345__24_), .Q(registers_a6_24_) );
	DFFPOSX1 DFFPOSX1_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17345__25_), .Q(registers_a6_25_) );
	DFFPOSX1 DFFPOSX1_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17345__26_), .Q(registers_a6_26_) );
	DFFPOSX1 DFFPOSX1_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17345__27_), .Q(registers_a6_27_) );
	DFFPOSX1 DFFPOSX1_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17345__28_), .Q(registers_a6_28_) );
	DFFPOSX1 DFFPOSX1_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17345__29_), .Q(registers_a6_29_) );
	DFFPOSX1 DFFPOSX1_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17345__30_), .Q(registers_a6_30_) );
	DFFPOSX1 DFFPOSX1_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17345__31_), .Q(registers_a6_31_) );
	DFFPOSX1 DFFPOSX1_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17346__0_), .Q(registers_a7_0_) );
	DFFPOSX1 DFFPOSX1_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17346__1_), .Q(registers_a7_1_) );
	DFFPOSX1 DFFPOSX1_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17346__2_), .Q(registers_a7_2_) );
	DFFPOSX1 DFFPOSX1_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17346__3_), .Q(registers_a7_3_) );
	DFFPOSX1 DFFPOSX1_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17346__4_), .Q(registers_a7_4_) );
	DFFPOSX1 DFFPOSX1_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17346__5_), .Q(registers_a7_5_) );
	DFFPOSX1 DFFPOSX1_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17346__6_), .Q(registers_a7_6_) );
	DFFPOSX1 DFFPOSX1_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17346__7_), .Q(registers_a7_7_) );
	DFFPOSX1 DFFPOSX1_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17346__8_), .Q(registers_a7_8_) );
	DFFPOSX1 DFFPOSX1_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17346__9_), .Q(registers_a7_9_) );
	DFFPOSX1 DFFPOSX1_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17346__10_), .Q(registers_a7_10_) );
	DFFPOSX1 DFFPOSX1_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17346__11_), .Q(registers_a7_11_) );
	DFFPOSX1 DFFPOSX1_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17346__12_), .Q(registers_a7_12_) );
	DFFPOSX1 DFFPOSX1_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17346__13_), .Q(registers_a7_13_) );
	DFFPOSX1 DFFPOSX1_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17346__14_), .Q(registers_a7_14_) );
	DFFPOSX1 DFFPOSX1_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17346__15_), .Q(registers_a7_15_) );
	DFFPOSX1 DFFPOSX1_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17346__16_), .Q(registers_a7_16_) );
	DFFPOSX1 DFFPOSX1_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17346__17_), .Q(registers_a7_17_) );
	DFFPOSX1 DFFPOSX1_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17346__18_), .Q(registers_a7_18_) );
	DFFPOSX1 DFFPOSX1_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17346__19_), .Q(registers_a7_19_) );
	DFFPOSX1 DFFPOSX1_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17346__20_), .Q(registers_a7_20_) );
	DFFPOSX1 DFFPOSX1_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17346__21_), .Q(registers_a7_21_) );
	DFFPOSX1 DFFPOSX1_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17346__22_), .Q(registers_a7_22_) );
	DFFPOSX1 DFFPOSX1_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17346__23_), .Q(registers_a7_23_) );
	DFFPOSX1 DFFPOSX1_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17346__24_), .Q(registers_a7_24_) );
	DFFPOSX1 DFFPOSX1_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17346__25_), .Q(registers_a7_25_) );
	DFFPOSX1 DFFPOSX1_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17346__26_), .Q(registers_a7_26_) );
	DFFPOSX1 DFFPOSX1_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17346__27_), .Q(registers_a7_27_) );
	DFFPOSX1 DFFPOSX1_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17346__28_), .Q(registers_a7_28_) );
	DFFPOSX1 DFFPOSX1_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17346__29_), .Q(registers_a7_29_) );
	DFFPOSX1 DFFPOSX1_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17346__30_), .Q(registers_a7_30_) );
	DFFPOSX1 DFFPOSX1_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17346__31_), .Q(registers_a7_31_) );
	DFFPOSX1 DFFPOSX1_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17347__0_), .Q(registers_r18_0_) );
	DFFPOSX1 DFFPOSX1_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17347__1_), .Q(registers_r18_1_) );
	DFFPOSX1 DFFPOSX1_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17347__2_), .Q(registers_r18_2_) );
	DFFPOSX1 DFFPOSX1_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17347__3_), .Q(registers_r18_3_) );
	DFFPOSX1 DFFPOSX1_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17347__4_), .Q(registers_r18_4_) );
	DFFPOSX1 DFFPOSX1_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17347__5_), .Q(registers_r18_5_) );
	DFFPOSX1 DFFPOSX1_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17347__6_), .Q(registers_r18_6_) );
	DFFPOSX1 DFFPOSX1_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17347__7_), .Q(registers_r18_7_) );
	DFFPOSX1 DFFPOSX1_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17347__8_), .Q(registers_r18_8_) );
	DFFPOSX1 DFFPOSX1_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17347__9_), .Q(registers_r18_9_) );
	DFFPOSX1 DFFPOSX1_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17347__10_), .Q(registers_r18_10_) );
	DFFPOSX1 DFFPOSX1_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17347__11_), .Q(registers_r18_11_) );
	DFFPOSX1 DFFPOSX1_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17347__12_), .Q(registers_r18_12_) );
	DFFPOSX1 DFFPOSX1_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17347__13_), .Q(registers_r18_13_) );
	DFFPOSX1 DFFPOSX1_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17347__14_), .Q(registers_r18_14_) );
	DFFPOSX1 DFFPOSX1_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17347__15_), .Q(registers_r18_15_) );
	DFFPOSX1 DFFPOSX1_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17347__16_), .Q(registers_r18_16_) );
	DFFPOSX1 DFFPOSX1_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17347__17_), .Q(registers_r18_17_) );
	DFFPOSX1 DFFPOSX1_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17347__18_), .Q(registers_r18_18_) );
	DFFPOSX1 DFFPOSX1_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17347__19_), .Q(registers_r18_19_) );
	DFFPOSX1 DFFPOSX1_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17347__20_), .Q(registers_r18_20_) );
	DFFPOSX1 DFFPOSX1_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17347__21_), .Q(registers_r18_21_) );
	DFFPOSX1 DFFPOSX1_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17347__22_), .Q(registers_r18_22_) );
	DFFPOSX1 DFFPOSX1_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17347__23_), .Q(registers_r18_23_) );
	DFFPOSX1 DFFPOSX1_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17347__24_), .Q(registers_r18_24_) );
	DFFPOSX1 DFFPOSX1_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17347__25_), .Q(registers_r18_25_) );
	DFFPOSX1 DFFPOSX1_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17347__26_), .Q(registers_r18_26_) );
	DFFPOSX1 DFFPOSX1_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17347__27_), .Q(registers_r18_27_) );
	DFFPOSX1 DFFPOSX1_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17347__28_), .Q(registers_r18_28_) );
	DFFPOSX1 DFFPOSX1_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17347__29_), .Q(registers_r18_29_) );
	DFFPOSX1 DFFPOSX1_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17347__30_), .Q(registers_r18_30_) );
	DFFPOSX1 DFFPOSX1_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17347__31_), .Q(registers_r18_31_) );
	DFFPOSX1 DFFPOSX1_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17348__0_), .Q(registers_r19_0_) );
	DFFPOSX1 DFFPOSX1_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17348__1_), .Q(registers_r19_1_) );
	DFFPOSX1 DFFPOSX1_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17348__2_), .Q(registers_r19_2_) );
	DFFPOSX1 DFFPOSX1_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17348__3_), .Q(registers_r19_3_) );
	DFFPOSX1 DFFPOSX1_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17348__4_), .Q(registers_r19_4_) );
	DFFPOSX1 DFFPOSX1_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17348__5_), .Q(registers_r19_5_) );
	DFFPOSX1 DFFPOSX1_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17348__6_), .Q(registers_r19_6_) );
	DFFPOSX1 DFFPOSX1_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17348__7_), .Q(registers_r19_7_) );
	DFFPOSX1 DFFPOSX1_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17348__8_), .Q(registers_r19_8_) );
	DFFPOSX1 DFFPOSX1_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17348__9_), .Q(registers_r19_9_) );
	DFFPOSX1 DFFPOSX1_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17348__10_), .Q(registers_r19_10_) );
	DFFPOSX1 DFFPOSX1_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17348__11_), .Q(registers_r19_11_) );
	DFFPOSX1 DFFPOSX1_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17348__12_), .Q(registers_r19_12_) );
	DFFPOSX1 DFFPOSX1_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17348__13_), .Q(registers_r19_13_) );
	DFFPOSX1 DFFPOSX1_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17348__14_), .Q(registers_r19_14_) );
	DFFPOSX1 DFFPOSX1_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17348__15_), .Q(registers_r19_15_) );
	DFFPOSX1 DFFPOSX1_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17348__16_), .Q(registers_r19_16_) );
	DFFPOSX1 DFFPOSX1_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17348__17_), .Q(registers_r19_17_) );
	DFFPOSX1 DFFPOSX1_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17348__18_), .Q(registers_r19_18_) );
	DFFPOSX1 DFFPOSX1_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17348__19_), .Q(registers_r19_19_) );
	DFFPOSX1 DFFPOSX1_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17348__20_), .Q(registers_r19_20_) );
	DFFPOSX1 DFFPOSX1_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17348__21_), .Q(registers_r19_21_) );
	DFFPOSX1 DFFPOSX1_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17348__22_), .Q(registers_r19_22_) );
	DFFPOSX1 DFFPOSX1_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17348__23_), .Q(registers_r19_23_) );
	DFFPOSX1 DFFPOSX1_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17348__24_), .Q(registers_r19_24_) );
	DFFPOSX1 DFFPOSX1_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17348__25_), .Q(registers_r19_25_) );
	DFFPOSX1 DFFPOSX1_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17348__26_), .Q(registers_r19_26_) );
	DFFPOSX1 DFFPOSX1_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17348__27_), .Q(registers_r19_27_) );
	DFFPOSX1 DFFPOSX1_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17348__28_), .Q(registers_r19_28_) );
	DFFPOSX1 DFFPOSX1_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17348__29_), .Q(registers_r19_29_) );
	DFFPOSX1 DFFPOSX1_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17348__30_), .Q(registers_r19_30_) );
	DFFPOSX1 DFFPOSX1_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17348__31_), .Q(registers_r19_31_) );
	DFFPOSX1 DFFPOSX1_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17350__0_), .Q(registers_r20_0_) );
	DFFPOSX1 DFFPOSX1_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17350__1_), .Q(registers_r20_1_) );
	DFFPOSX1 DFFPOSX1_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17350__2_), .Q(registers_r20_2_) );
	DFFPOSX1 DFFPOSX1_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17350__3_), .Q(registers_r20_3_) );
	DFFPOSX1 DFFPOSX1_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17350__4_), .Q(registers_r20_4_) );
	DFFPOSX1 DFFPOSX1_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17350__5_), .Q(registers_r20_5_) );
	DFFPOSX1 DFFPOSX1_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17350__6_), .Q(registers_r20_6_) );
	DFFPOSX1 DFFPOSX1_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17350__7_), .Q(registers_r20_7_) );
	DFFPOSX1 DFFPOSX1_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17350__8_), .Q(registers_r20_8_) );
	DFFPOSX1 DFFPOSX1_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17350__9_), .Q(registers_r20_9_) );
	DFFPOSX1 DFFPOSX1_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17350__10_), .Q(registers_r20_10_) );
	DFFPOSX1 DFFPOSX1_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17350__11_), .Q(registers_r20_11_) );
	DFFPOSX1 DFFPOSX1_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17350__12_), .Q(registers_r20_12_) );
	DFFPOSX1 DFFPOSX1_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17350__13_), .Q(registers_r20_13_) );
	DFFPOSX1 DFFPOSX1_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17350__14_), .Q(registers_r20_14_) );
	DFFPOSX1 DFFPOSX1_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17350__15_), .Q(registers_r20_15_) );
	DFFPOSX1 DFFPOSX1_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17350__16_), .Q(registers_r20_16_) );
	DFFPOSX1 DFFPOSX1_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17350__17_), .Q(registers_r20_17_) );
	DFFPOSX1 DFFPOSX1_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17350__18_), .Q(registers_r20_18_) );
	DFFPOSX1 DFFPOSX1_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17350__19_), .Q(registers_r20_19_) );
	DFFPOSX1 DFFPOSX1_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17350__20_), .Q(registers_r20_20_) );
	DFFPOSX1 DFFPOSX1_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17350__21_), .Q(registers_r20_21_) );
	DFFPOSX1 DFFPOSX1_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17350__22_), .Q(registers_r20_22_) );
	DFFPOSX1 DFFPOSX1_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17350__23_), .Q(registers_r20_23_) );
	DFFPOSX1 DFFPOSX1_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17350__24_), .Q(registers_r20_24_) );
	DFFPOSX1 DFFPOSX1_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17350__25_), .Q(registers_r20_25_) );
	DFFPOSX1 DFFPOSX1_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17350__26_), .Q(registers_r20_26_) );
	DFFPOSX1 DFFPOSX1_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17350__27_), .Q(registers_r20_27_) );
	DFFPOSX1 DFFPOSX1_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17350__28_), .Q(registers_r20_28_) );
	DFFPOSX1 DFFPOSX1_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17350__29_), .Q(registers_r20_29_) );
	DFFPOSX1 DFFPOSX1_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17350__30_), .Q(registers_r20_30_) );
	DFFPOSX1 DFFPOSX1_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17350__31_), .Q(registers_r20_31_) );
	DFFPOSX1 DFFPOSX1_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17351__0_), .Q(registers_r21_0_) );
	DFFPOSX1 DFFPOSX1_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17351__1_), .Q(registers_r21_1_) );
	DFFPOSX1 DFFPOSX1_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17351__2_), .Q(registers_r21_2_) );
	DFFPOSX1 DFFPOSX1_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17351__3_), .Q(registers_r21_3_) );
	DFFPOSX1 DFFPOSX1_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17351__4_), .Q(registers_r21_4_) );
	DFFPOSX1 DFFPOSX1_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17351__5_), .Q(registers_r21_5_) );
	DFFPOSX1 DFFPOSX1_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17351__6_), .Q(registers_r21_6_) );
	DFFPOSX1 DFFPOSX1_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17351__7_), .Q(registers_r21_7_) );
	DFFPOSX1 DFFPOSX1_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17351__8_), .Q(registers_r21_8_) );
	DFFPOSX1 DFFPOSX1_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17351__9_), .Q(registers_r21_9_) );
	DFFPOSX1 DFFPOSX1_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17351__10_), .Q(registers_r21_10_) );
	DFFPOSX1 DFFPOSX1_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17351__11_), .Q(registers_r21_11_) );
	DFFPOSX1 DFFPOSX1_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17351__12_), .Q(registers_r21_12_) );
	DFFPOSX1 DFFPOSX1_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17351__13_), .Q(registers_r21_13_) );
	DFFPOSX1 DFFPOSX1_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17351__14_), .Q(registers_r21_14_) );
	DFFPOSX1 DFFPOSX1_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17351__15_), .Q(registers_r21_15_) );
	DFFPOSX1 DFFPOSX1_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17351__16_), .Q(registers_r21_16_) );
	DFFPOSX1 DFFPOSX1_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17351__17_), .Q(registers_r21_17_) );
	DFFPOSX1 DFFPOSX1_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17351__18_), .Q(registers_r21_18_) );
	DFFPOSX1 DFFPOSX1_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17351__19_), .Q(registers_r21_19_) );
	DFFPOSX1 DFFPOSX1_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17351__20_), .Q(registers_r21_20_) );
	DFFPOSX1 DFFPOSX1_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17351__21_), .Q(registers_r21_21_) );
	DFFPOSX1 DFFPOSX1_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17351__22_), .Q(registers_r21_22_) );
	DFFPOSX1 DFFPOSX1_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17351__23_), .Q(registers_r21_23_) );
	DFFPOSX1 DFFPOSX1_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17351__24_), .Q(registers_r21_24_) );
	DFFPOSX1 DFFPOSX1_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17351__25_), .Q(registers_r21_25_) );
	DFFPOSX1 DFFPOSX1_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17351__26_), .Q(registers_r21_26_) );
	DFFPOSX1 DFFPOSX1_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17351__27_), .Q(registers_r21_27_) );
	DFFPOSX1 DFFPOSX1_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17351__28_), .Q(registers_r21_28_) );
	DFFPOSX1 DFFPOSX1_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17351__29_), .Q(registers_r21_29_) );
	DFFPOSX1 DFFPOSX1_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17351__30_), .Q(registers_r21_30_) );
	DFFPOSX1 DFFPOSX1_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17351__31_), .Q(registers_r21_31_) );
	DFFPOSX1 DFFPOSX1_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17352__0_), .Q(registers_r22_0_) );
	DFFPOSX1 DFFPOSX1_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17352__1_), .Q(registers_r22_1_) );
	DFFPOSX1 DFFPOSX1_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17352__2_), .Q(registers_r22_2_) );
	DFFPOSX1 DFFPOSX1_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17352__3_), .Q(registers_r22_3_) );
	DFFPOSX1 DFFPOSX1_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17352__4_), .Q(registers_r22_4_) );
	DFFPOSX1 DFFPOSX1_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17352__5_), .Q(registers_r22_5_) );
	DFFPOSX1 DFFPOSX1_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17352__6_), .Q(registers_r22_6_) );
	DFFPOSX1 DFFPOSX1_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17352__7_), .Q(registers_r22_7_) );
	DFFPOSX1 DFFPOSX1_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17352__8_), .Q(registers_r22_8_) );
	DFFPOSX1 DFFPOSX1_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17352__9_), .Q(registers_r22_9_) );
	DFFPOSX1 DFFPOSX1_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17352__10_), .Q(registers_r22_10_) );
	DFFPOSX1 DFFPOSX1_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17352__11_), .Q(registers_r22_11_) );
	DFFPOSX1 DFFPOSX1_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17352__12_), .Q(registers_r22_12_) );
	DFFPOSX1 DFFPOSX1_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17352__13_), .Q(registers_r22_13_) );
	DFFPOSX1 DFFPOSX1_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17352__14_), .Q(registers_r22_14_) );
	DFFPOSX1 DFFPOSX1_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17352__15_), .Q(registers_r22_15_) );
	DFFPOSX1 DFFPOSX1_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17352__16_), .Q(registers_r22_16_) );
	DFFPOSX1 DFFPOSX1_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17352__17_), .Q(registers_r22_17_) );
	DFFPOSX1 DFFPOSX1_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17352__18_), .Q(registers_r22_18_) );
	DFFPOSX1 DFFPOSX1_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17352__19_), .Q(registers_r22_19_) );
	DFFPOSX1 DFFPOSX1_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17352__20_), .Q(registers_r22_20_) );
	DFFPOSX1 DFFPOSX1_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17352__21_), .Q(registers_r22_21_) );
	DFFPOSX1 DFFPOSX1_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17352__22_), .Q(registers_r22_22_) );
	DFFPOSX1 DFFPOSX1_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17352__23_), .Q(registers_r22_23_) );
	DFFPOSX1 DFFPOSX1_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17352__24_), .Q(registers_r22_24_) );
	DFFPOSX1 DFFPOSX1_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17352__25_), .Q(registers_r22_25_) );
	DFFPOSX1 DFFPOSX1_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17352__26_), .Q(registers_r22_26_) );
	DFFPOSX1 DFFPOSX1_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17352__27_), .Q(registers_r22_27_) );
	DFFPOSX1 DFFPOSX1_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17352__28_), .Q(registers_r22_28_) );
	DFFPOSX1 DFFPOSX1_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17352__29_), .Q(registers_r22_29_) );
	DFFPOSX1 DFFPOSX1_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17352__30_), .Q(registers_r22_30_) );
	DFFPOSX1 DFFPOSX1_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17352__31_), .Q(registers_r22_31_) );
	DFFPOSX1 DFFPOSX1_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17353__0_), .Q(registers_r23_0_) );
	DFFPOSX1 DFFPOSX1_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17353__1_), .Q(registers_r23_1_) );
	DFFPOSX1 DFFPOSX1_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17353__2_), .Q(registers_r23_2_) );
	DFFPOSX1 DFFPOSX1_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17353__3_), .Q(registers_r23_3_) );
	DFFPOSX1 DFFPOSX1_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17353__4_), .Q(registers_r23_4_) );
	DFFPOSX1 DFFPOSX1_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17353__5_), .Q(registers_r23_5_) );
	DFFPOSX1 DFFPOSX1_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17353__6_), .Q(registers_r23_6_) );
	DFFPOSX1 DFFPOSX1_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17353__7_), .Q(registers_r23_7_) );
	DFFPOSX1 DFFPOSX1_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17353__8_), .Q(registers_r23_8_) );
	DFFPOSX1 DFFPOSX1_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17353__9_), .Q(registers_r23_9_) );
	DFFPOSX1 DFFPOSX1_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17353__10_), .Q(registers_r23_10_) );
	DFFPOSX1 DFFPOSX1_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17353__11_), .Q(registers_r23_11_) );
	DFFPOSX1 DFFPOSX1_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17353__12_), .Q(registers_r23_12_) );
	DFFPOSX1 DFFPOSX1_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17353__13_), .Q(registers_r23_13_) );
	DFFPOSX1 DFFPOSX1_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17353__14_), .Q(registers_r23_14_) );
	DFFPOSX1 DFFPOSX1_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17353__15_), .Q(registers_r23_15_) );
	DFFPOSX1 DFFPOSX1_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17353__16_), .Q(registers_r23_16_) );
	DFFPOSX1 DFFPOSX1_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17353__17_), .Q(registers_r23_17_) );
	DFFPOSX1 DFFPOSX1_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17353__18_), .Q(registers_r23_18_) );
	DFFPOSX1 DFFPOSX1_845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17353__19_), .Q(registers_r23_19_) );
	DFFPOSX1 DFFPOSX1_846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17353__20_), .Q(registers_r23_20_) );
	DFFPOSX1 DFFPOSX1_847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17353__21_), .Q(registers_r23_21_) );
	DFFPOSX1 DFFPOSX1_848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17353__22_), .Q(registers_r23_22_) );
	DFFPOSX1 DFFPOSX1_849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17353__23_), .Q(registers_r23_23_) );
	DFFPOSX1 DFFPOSX1_850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17353__24_), .Q(registers_r23_24_) );
	DFFPOSX1 DFFPOSX1_851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17353__25_), .Q(registers_r23_25_) );
	DFFPOSX1 DFFPOSX1_852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17353__26_), .Q(registers_r23_26_) );
	DFFPOSX1 DFFPOSX1_853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17353__27_), .Q(registers_r23_27_) );
	DFFPOSX1 DFFPOSX1_854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17353__28_), .Q(registers_r23_28_) );
	DFFPOSX1 DFFPOSX1_855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17353__29_), .Q(registers_r23_29_) );
	DFFPOSX1 DFFPOSX1_856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17353__30_), .Q(registers_r23_30_) );
	DFFPOSX1 DFFPOSX1_857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17353__31_), .Q(registers_r23_31_) );
	DFFPOSX1 DFFPOSX1_858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17354__0_), .Q(registers_r24_0_) );
	DFFPOSX1 DFFPOSX1_859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17354__1_), .Q(registers_r24_1_) );
	DFFPOSX1 DFFPOSX1_860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17354__2_), .Q(registers_r24_2_) );
	DFFPOSX1 DFFPOSX1_861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17354__3_), .Q(registers_r24_3_) );
	DFFPOSX1 DFFPOSX1_862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17354__4_), .Q(registers_r24_4_) );
	DFFPOSX1 DFFPOSX1_863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17354__5_), .Q(registers_r24_5_) );
	DFFPOSX1 DFFPOSX1_864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17354__6_), .Q(registers_r24_6_) );
	DFFPOSX1 DFFPOSX1_865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17354__7_), .Q(registers_r24_7_) );
	DFFPOSX1 DFFPOSX1_866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17354__8_), .Q(registers_r24_8_) );
	DFFPOSX1 DFFPOSX1_867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17354__9_), .Q(registers_r24_9_) );
	DFFPOSX1 DFFPOSX1_868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17354__10_), .Q(registers_r24_10_) );
	DFFPOSX1 DFFPOSX1_869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17354__11_), .Q(registers_r24_11_) );
	DFFPOSX1 DFFPOSX1_870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17354__12_), .Q(registers_r24_12_) );
	DFFPOSX1 DFFPOSX1_871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17354__13_), .Q(registers_r24_13_) );
	DFFPOSX1 DFFPOSX1_872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17354__14_), .Q(registers_r24_14_) );
	DFFPOSX1 DFFPOSX1_873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17354__15_), .Q(registers_r24_15_) );
	DFFPOSX1 DFFPOSX1_874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17354__16_), .Q(registers_r24_16_) );
	DFFPOSX1 DFFPOSX1_875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17354__17_), .Q(registers_r24_17_) );
	DFFPOSX1 DFFPOSX1_876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17354__18_), .Q(registers_r24_18_) );
	DFFPOSX1 DFFPOSX1_877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17354__19_), .Q(registers_r24_19_) );
	DFFPOSX1 DFFPOSX1_878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17354__20_), .Q(registers_r24_20_) );
	DFFPOSX1 DFFPOSX1_879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17354__21_), .Q(registers_r24_21_) );
	DFFPOSX1 DFFPOSX1_880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17354__22_), .Q(registers_r24_22_) );
	DFFPOSX1 DFFPOSX1_881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17354__23_), .Q(registers_r24_23_) );
	DFFPOSX1 DFFPOSX1_882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17354__24_), .Q(registers_r24_24_) );
	DFFPOSX1 DFFPOSX1_883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17354__25_), .Q(registers_r24_25_) );
	DFFPOSX1 DFFPOSX1_884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17354__26_), .Q(registers_r24_26_) );
	DFFPOSX1 DFFPOSX1_885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17354__27_), .Q(registers_r24_27_) );
	DFFPOSX1 DFFPOSX1_886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17354__28_), .Q(registers_r24_28_) );
	DFFPOSX1 DFFPOSX1_887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17354__29_), .Q(registers_r24_29_) );
	DFFPOSX1 DFFPOSX1_888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17354__30_), .Q(registers_r24_30_) );
	DFFPOSX1 DFFPOSX1_889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17354__31_), .Q(registers_r24_31_) );
	DFFPOSX1 DFFPOSX1_890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17355__0_), .Q(registers_r25_0_) );
	DFFPOSX1 DFFPOSX1_891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17355__1_), .Q(registers_r25_1_) );
	DFFPOSX1 DFFPOSX1_892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17355__2_), .Q(registers_r25_2_) );
	DFFPOSX1 DFFPOSX1_893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17355__3_), .Q(registers_r25_3_) );
	DFFPOSX1 DFFPOSX1_894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17355__4_), .Q(registers_r25_4_) );
	DFFPOSX1 DFFPOSX1_895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17355__5_), .Q(registers_r25_5_) );
	DFFPOSX1 DFFPOSX1_896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17355__6_), .Q(registers_r25_6_) );
	DFFPOSX1 DFFPOSX1_897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17355__7_), .Q(registers_r25_7_) );
	DFFPOSX1 DFFPOSX1_898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17355__8_), .Q(registers_r25_8_) );
	DFFPOSX1 DFFPOSX1_899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17355__9_), .Q(registers_r25_9_) );
	DFFPOSX1 DFFPOSX1_900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17355__10_), .Q(registers_r25_10_) );
	DFFPOSX1 DFFPOSX1_901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17355__11_), .Q(registers_r25_11_) );
	DFFPOSX1 DFFPOSX1_902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17355__12_), .Q(registers_r25_12_) );
	DFFPOSX1 DFFPOSX1_903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17355__13_), .Q(registers_r25_13_) );
	DFFPOSX1 DFFPOSX1_904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17355__14_), .Q(registers_r25_14_) );
	DFFPOSX1 DFFPOSX1_905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17355__15_), .Q(registers_r25_15_) );
	DFFPOSX1 DFFPOSX1_906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17355__16_), .Q(registers_r25_16_) );
	DFFPOSX1 DFFPOSX1_907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17355__17_), .Q(registers_r25_17_) );
	DFFPOSX1 DFFPOSX1_908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17355__18_), .Q(registers_r25_18_) );
	DFFPOSX1 DFFPOSX1_909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17355__19_), .Q(registers_r25_19_) );
	DFFPOSX1 DFFPOSX1_910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17355__20_), .Q(registers_r25_20_) );
	DFFPOSX1 DFFPOSX1_911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17355__21_), .Q(registers_r25_21_) );
	DFFPOSX1 DFFPOSX1_912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17355__22_), .Q(registers_r25_22_) );
	DFFPOSX1 DFFPOSX1_913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17355__23_), .Q(registers_r25_23_) );
	DFFPOSX1 DFFPOSX1_914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17355__24_), .Q(registers_r25_24_) );
	DFFPOSX1 DFFPOSX1_915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17355__25_), .Q(registers_r25_25_) );
	DFFPOSX1 DFFPOSX1_916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17355__26_), .Q(registers_r25_26_) );
	DFFPOSX1 DFFPOSX1_917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17355__27_), .Q(registers_r25_27_) );
	DFFPOSX1 DFFPOSX1_918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17355__28_), .Q(registers_r25_28_) );
	DFFPOSX1 DFFPOSX1_919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17355__29_), .Q(registers_r25_29_) );
	DFFPOSX1 DFFPOSX1_920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17355__30_), .Q(registers_r25_30_) );
	DFFPOSX1 DFFPOSX1_921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17355__31_), .Q(registers_r25_31_) );
	DFFPOSX1 DFFPOSX1_922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17356__0_), .Q(registers_r26_0_) );
	DFFPOSX1 DFFPOSX1_923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17356__1_), .Q(registers_r26_1_) );
	DFFPOSX1 DFFPOSX1_924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17356__2_), .Q(registers_r26_2_) );
	DFFPOSX1 DFFPOSX1_925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17356__3_), .Q(registers_r26_3_) );
	DFFPOSX1 DFFPOSX1_926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17356__4_), .Q(registers_r26_4_) );
	DFFPOSX1 DFFPOSX1_927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17356__5_), .Q(registers_r26_5_) );
	DFFPOSX1 DFFPOSX1_928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17356__6_), .Q(registers_r26_6_) );
	DFFPOSX1 DFFPOSX1_929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17356__7_), .Q(registers_r26_7_) );
	DFFPOSX1 DFFPOSX1_930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17356__8_), .Q(registers_r26_8_) );
	DFFPOSX1 DFFPOSX1_931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17356__9_), .Q(registers_r26_9_) );
	DFFPOSX1 DFFPOSX1_932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17356__10_), .Q(registers_r26_10_) );
	DFFPOSX1 DFFPOSX1_933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17356__11_), .Q(registers_r26_11_) );
	DFFPOSX1 DFFPOSX1_934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17356__12_), .Q(registers_r26_12_) );
	DFFPOSX1 DFFPOSX1_935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17356__13_), .Q(registers_r26_13_) );
	DFFPOSX1 DFFPOSX1_936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17356__14_), .Q(registers_r26_14_) );
	DFFPOSX1 DFFPOSX1_937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17356__15_), .Q(registers_r26_15_) );
	DFFPOSX1 DFFPOSX1_938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17356__16_), .Q(registers_r26_16_) );
	DFFPOSX1 DFFPOSX1_939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17356__17_), .Q(registers_r26_17_) );
	DFFPOSX1 DFFPOSX1_940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17356__18_), .Q(registers_r26_18_) );
	DFFPOSX1 DFFPOSX1_941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17356__19_), .Q(registers_r26_19_) );
	DFFPOSX1 DFFPOSX1_942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17356__20_), .Q(registers_r26_20_) );
	DFFPOSX1 DFFPOSX1_943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17356__21_), .Q(registers_r26_21_) );
	DFFPOSX1 DFFPOSX1_944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17356__22_), .Q(registers_r26_22_) );
	DFFPOSX1 DFFPOSX1_945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17356__23_), .Q(registers_r26_23_) );
	DFFPOSX1 DFFPOSX1_946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17356__24_), .Q(registers_r26_24_) );
	DFFPOSX1 DFFPOSX1_947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17356__25_), .Q(registers_r26_25_) );
	DFFPOSX1 DFFPOSX1_948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17356__26_), .Q(registers_r26_26_) );
	DFFPOSX1 DFFPOSX1_949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17356__27_), .Q(registers_r26_27_) );
	DFFPOSX1 DFFPOSX1_950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17356__28_), .Q(registers_r26_28_) );
	DFFPOSX1 DFFPOSX1_951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17356__29_), .Q(registers_r26_29_) );
	DFFPOSX1 DFFPOSX1_952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17356__30_), .Q(registers_r26_30_) );
	DFFPOSX1 DFFPOSX1_953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17356__31_), .Q(registers_r26_31_) );
	DFFPOSX1 DFFPOSX1_954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17357__0_), .Q(registers_r27_0_) );
	DFFPOSX1 DFFPOSX1_955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17357__1_), .Q(registers_r27_1_) );
	DFFPOSX1 DFFPOSX1_956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17357__2_), .Q(registers_r27_2_) );
	DFFPOSX1 DFFPOSX1_957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17357__3_), .Q(registers_r27_3_) );
	DFFPOSX1 DFFPOSX1_958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17357__4_), .Q(registers_r27_4_) );
	DFFPOSX1 DFFPOSX1_959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17357__5_), .Q(registers_r27_5_) );
	DFFPOSX1 DFFPOSX1_960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17357__6_), .Q(registers_r27_6_) );
	DFFPOSX1 DFFPOSX1_961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17357__7_), .Q(registers_r27_7_) );
	DFFPOSX1 DFFPOSX1_962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17357__8_), .Q(registers_r27_8_) );
	DFFPOSX1 DFFPOSX1_963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17357__9_), .Q(registers_r27_9_) );
	DFFPOSX1 DFFPOSX1_964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17357__10_), .Q(registers_r27_10_) );
	DFFPOSX1 DFFPOSX1_965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17357__11_), .Q(registers_r27_11_) );
	DFFPOSX1 DFFPOSX1_966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17357__12_), .Q(registers_r27_12_) );
	DFFPOSX1 DFFPOSX1_967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17357__13_), .Q(registers_r27_13_) );
	DFFPOSX1 DFFPOSX1_968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17357__14_), .Q(registers_r27_14_) );
	DFFPOSX1 DFFPOSX1_969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17357__15_), .Q(registers_r27_15_) );
	DFFPOSX1 DFFPOSX1_970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17357__16_), .Q(registers_r27_16_) );
	DFFPOSX1 DFFPOSX1_971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17357__17_), .Q(registers_r27_17_) );
	DFFPOSX1 DFFPOSX1_972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17357__18_), .Q(registers_r27_18_) );
	DFFPOSX1 DFFPOSX1_973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17357__19_), .Q(registers_r27_19_) );
	DFFPOSX1 DFFPOSX1_974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17357__20_), .Q(registers_r27_20_) );
	DFFPOSX1 DFFPOSX1_975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17357__21_), .Q(registers_r27_21_) );
	DFFPOSX1 DFFPOSX1_976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17357__22_), .Q(registers_r27_22_) );
	DFFPOSX1 DFFPOSX1_977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17357__23_), .Q(registers_r27_23_) );
	DFFPOSX1 DFFPOSX1_978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17357__24_), .Q(registers_r27_24_) );
	DFFPOSX1 DFFPOSX1_979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17357__25_), .Q(registers_r27_25_) );
	DFFPOSX1 DFFPOSX1_980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17357__26_), .Q(registers_r27_26_) );
	DFFPOSX1 DFFPOSX1_981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17357__27_), .Q(registers_r27_27_) );
	DFFPOSX1 DFFPOSX1_982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17357__28_), .Q(registers_r27_28_) );
	DFFPOSX1 DFFPOSX1_983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17357__29_), .Q(registers_r27_29_) );
	DFFPOSX1 DFFPOSX1_984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17357__30_), .Q(registers_r27_30_) );
	DFFPOSX1 DFFPOSX1_985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17357__31_), .Q(registers_r27_31_) );
	DFFPOSX1 DFFPOSX1_986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17358__0_), .Q(registers_r28_0_) );
	DFFPOSX1 DFFPOSX1_987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17358__1_), .Q(registers_r28_1_) );
	DFFPOSX1 DFFPOSX1_988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17358__2_), .Q(registers_r28_2_) );
	DFFPOSX1 DFFPOSX1_989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17358__3_), .Q(registers_r28_3_) );
	DFFPOSX1 DFFPOSX1_990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17358__4_), .Q(registers_r28_4_) );
	DFFPOSX1 DFFPOSX1_991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17358__5_), .Q(registers_r28_5_) );
	DFFPOSX1 DFFPOSX1_992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17358__6_), .Q(registers_r28_6_) );
	DFFPOSX1 DFFPOSX1_993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17358__7_), .Q(registers_r28_7_) );
	DFFPOSX1 DFFPOSX1_994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17358__8_), .Q(registers_r28_8_) );
	DFFPOSX1 DFFPOSX1_995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17358__9_), .Q(registers_r28_9_) );
	DFFPOSX1 DFFPOSX1_996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17358__10_), .Q(registers_r28_10_) );
	DFFPOSX1 DFFPOSX1_997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17358__11_), .Q(registers_r28_11_) );
	DFFPOSX1 DFFPOSX1_998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17358__12_), .Q(registers_r28_12_) );
	DFFPOSX1 DFFPOSX1_999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17358__13_), .Q(registers_r28_13_) );
	DFFPOSX1 DFFPOSX1_1000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17358__14_), .Q(registers_r28_14_) );
	DFFPOSX1 DFFPOSX1_1001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17358__15_), .Q(registers_r28_15_) );
	DFFPOSX1 DFFPOSX1_1002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17358__16_), .Q(registers_r28_16_) );
	DFFPOSX1 DFFPOSX1_1003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17358__17_), .Q(registers_r28_17_) );
	DFFPOSX1 DFFPOSX1_1004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17358__18_), .Q(registers_r28_18_) );
	DFFPOSX1 DFFPOSX1_1005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17358__19_), .Q(registers_r28_19_) );
	DFFPOSX1 DFFPOSX1_1006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17358__20_), .Q(registers_r28_20_) );
	DFFPOSX1 DFFPOSX1_1007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_17358__21_), .Q(registers_r28_21_) );
	DFFPOSX1 DFFPOSX1_1008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_17358__22_), .Q(registers_r28_22_) );
	DFFPOSX1 DFFPOSX1_1009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_17358__23_), .Q(registers_r28_23_) );
	DFFPOSX1 DFFPOSX1_1010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_17358__24_), .Q(registers_r28_24_) );
	DFFPOSX1 DFFPOSX1_1011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_17358__25_), .Q(registers_r28_25_) );
	DFFPOSX1 DFFPOSX1_1012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_17358__26_), .Q(registers_r28_26_) );
	DFFPOSX1 DFFPOSX1_1013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_17358__27_), .Q(registers_r28_27_) );
	DFFPOSX1 DFFPOSX1_1014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_17358__28_), .Q(registers_r28_28_) );
	DFFPOSX1 DFFPOSX1_1015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_17358__29_), .Q(registers_r28_29_) );
	DFFPOSX1 DFFPOSX1_1016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_17358__30_), .Q(registers_r28_30_) );
	DFFPOSX1 DFFPOSX1_1017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_17358__31_), .Q(registers_r28_31_) );
	DFFPOSX1 DFFPOSX1_1018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_17359__0_), .Q(registers_r29_0_) );
	DFFPOSX1 DFFPOSX1_1019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_17359__1_), .Q(registers_r29_1_) );
	DFFPOSX1 DFFPOSX1_1020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_17359__2_), .Q(registers_r29_2_) );
	DFFPOSX1 DFFPOSX1_1021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_17359__3_), .Q(registers_r29_3_) );
	DFFPOSX1 DFFPOSX1_1022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_17359__4_), .Q(registers_r29_4_) );
	DFFPOSX1 DFFPOSX1_1023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_17359__5_), .Q(registers_r29_5_) );
	DFFPOSX1 DFFPOSX1_1024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_17359__6_), .Q(registers_r29_6_) );
	DFFPOSX1 DFFPOSX1_1025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_17359__7_), .Q(registers_r29_7_) );
	DFFPOSX1 DFFPOSX1_1026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_17359__8_), .Q(registers_r29_8_) );
	DFFPOSX1 DFFPOSX1_1027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_17359__9_), .Q(registers_r29_9_) );
	DFFPOSX1 DFFPOSX1_1028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_17359__10_), .Q(registers_r29_10_) );
	DFFPOSX1 DFFPOSX1_1029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17359__11_), .Q(registers_r29_11_) );
	DFFPOSX1 DFFPOSX1_1030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_17359__12_), .Q(registers_r29_12_) );
	DFFPOSX1 DFFPOSX1_1031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17359__13_), .Q(registers_r29_13_) );
	DFFPOSX1 DFFPOSX1_1032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_17359__14_), .Q(registers_r29_14_) );
	DFFPOSX1 DFFPOSX1_1033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_17359__15_), .Q(registers_r29_15_) );
	DFFPOSX1 DFFPOSX1_1034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_17359__16_), .Q(registers_r29_16_) );
	DFFPOSX1 DFFPOSX1_1035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_17359__17_), .Q(registers_r29_17_) );
	DFFPOSX1 DFFPOSX1_1036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_17359__18_), .Q(registers_r29_18_) );
	DFFPOSX1 DFFPOSX1_1037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_17359__19_), .Q(registers_r29_19_) );
	DFFPOSX1 DFFPOSX1_1038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_17359__20_), .Q(registers_r29_20_) );
	DFFPOSX1 DFFPOSX1_1039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_17359__21_), .Q(registers_r29_21_) );
	DFFPOSX1 DFFPOSX1_1040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_17359__22_), .Q(registers_r29_22_) );
	DFFPOSX1 DFFPOSX1_1041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_17359__23_), .Q(registers_r29_23_) );
	DFFPOSX1 DFFPOSX1_1042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_17359__24_), .Q(registers_r29_24_) );
	DFFPOSX1 DFFPOSX1_1043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_17359__25_), .Q(registers_r29_25_) );
	DFFPOSX1 DFFPOSX1_1044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_17359__26_), .Q(registers_r29_26_) );
	DFFPOSX1 DFFPOSX1_1045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_17359__27_), .Q(registers_r29_27_) );
	DFFPOSX1 DFFPOSX1_1046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_17359__28_), .Q(registers_r29_28_) );
	DFFPOSX1 DFFPOSX1_1047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_17359__29_), .Q(registers_r29_29_) );
	DFFPOSX1 DFFPOSX1_1048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_17359__30_), .Q(registers_r29_30_) );
	DFFPOSX1 DFFPOSX1_1049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_17359__31_), .Q(registers_r29_31_) );
	DFFPOSX1 DFFPOSX1_1050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_17361__0_), .Q(registers_r30_0_) );
	DFFPOSX1 DFFPOSX1_1051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_17361__1_), .Q(registers_r30_1_) );
	DFFPOSX1 DFFPOSX1_1052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_17361__2_), .Q(registers_r30_2_) );
	DFFPOSX1 DFFPOSX1_1053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_17361__3_), .Q(registers_r30_3_) );
	DFFPOSX1 DFFPOSX1_1054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_17361__4_), .Q(registers_r30_4_) );
	DFFPOSX1 DFFPOSX1_1055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_17361__5_), .Q(registers_r30_5_) );
	DFFPOSX1 DFFPOSX1_1056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_17361__6_), .Q(registers_r30_6_) );
	DFFPOSX1 DFFPOSX1_1057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_17361__7_), .Q(registers_r30_7_) );
	DFFPOSX1 DFFPOSX1_1058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_17361__8_), .Q(registers_r30_8_) );
	DFFPOSX1 DFFPOSX1_1059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_17361__9_), .Q(registers_r30_9_) );
	DFFPOSX1 DFFPOSX1_1060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_17361__10_), .Q(registers_r30_10_) );
	DFFPOSX1 DFFPOSX1_1061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_17361__11_), .Q(registers_r30_11_) );
	DFFPOSX1 DFFPOSX1_1062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_17361__12_), .Q(registers_r30_12_) );
	DFFPOSX1 DFFPOSX1_1063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_17361__13_), .Q(registers_r30_13_) );
	DFFPOSX1 DFFPOSX1_1064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_17361__14_), .Q(registers_r30_14_) );
	DFFPOSX1 DFFPOSX1_1065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_17361__15_), .Q(registers_r30_15_) );
	DFFPOSX1 DFFPOSX1_1066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_17361__16_), .Q(registers_r30_16_) );
	DFFPOSX1 DFFPOSX1_1067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17361__17_), .Q(registers_r30_17_) );
	DFFPOSX1 DFFPOSX1_1068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_17361__18_), .Q(registers_r30_18_) );
	DFFPOSX1 DFFPOSX1_1069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_17361__19_), .Q(registers_r30_19_) );
	DFFPOSX1 DFFPOSX1_1070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_17361__20_), .Q(registers_r30_20_) );
	DFFPOSX1 DFFPOSX1_1071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_17361__21_), .Q(registers_r30_21_) );
	DFFPOSX1 DFFPOSX1_1072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_17361__22_), .Q(registers_r30_22_) );
	DFFPOSX1 DFFPOSX1_1073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_17361__23_), .Q(registers_r30_23_) );
	DFFPOSX1 DFFPOSX1_1074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_17361__24_), .Q(registers_r30_24_) );
	DFFPOSX1 DFFPOSX1_1075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_17361__25_), .Q(registers_r30_25_) );
	DFFPOSX1 DFFPOSX1_1076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_17361__26_), .Q(registers_r30_26_) );
	DFFPOSX1 DFFPOSX1_1077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_17361__27_), .Q(registers_r30_27_) );
	DFFPOSX1 DFFPOSX1_1078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_17361__28_), .Q(registers_r30_28_) );
	DFFPOSX1 DFFPOSX1_1079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_17361__29_), .Q(registers_r30_29_) );
	DFFPOSX1 DFFPOSX1_1080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_17361__30_), .Q(registers_r30_30_) );
	DFFPOSX1 DFFPOSX1_1081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_17361__31_), .Q(registers_r30_31_) );
	DFFPOSX1 DFFPOSX1_1082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_17362__0_), .Q(registers_r31_0_) );
	DFFPOSX1 DFFPOSX1_1083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_17362__1_), .Q(registers_r31_1_) );
	DFFPOSX1 DFFPOSX1_1084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_17362__2_), .Q(registers_r31_2_) );
	DFFPOSX1 DFFPOSX1_1085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_17362__3_), .Q(registers_r31_3_) );
	DFFPOSX1 DFFPOSX1_1086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_17362__4_), .Q(registers_r31_4_) );
	DFFPOSX1 DFFPOSX1_1087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_17362__5_), .Q(registers_r31_5_) );
	DFFPOSX1 DFFPOSX1_1088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_17362__6_), .Q(registers_r31_6_) );
	DFFPOSX1 DFFPOSX1_1089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_17362__7_), .Q(registers_r31_7_) );
	DFFPOSX1 DFFPOSX1_1090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_17362__8_), .Q(registers_r31_8_) );
	DFFPOSX1 DFFPOSX1_1091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_17362__9_), .Q(registers_r31_9_) );
	DFFPOSX1 DFFPOSX1_1092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_17362__10_), .Q(registers_r31_10_) );
	DFFPOSX1 DFFPOSX1_1093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_17362__11_), .Q(registers_r31_11_) );
	DFFPOSX1 DFFPOSX1_1094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_17362__12_), .Q(registers_r31_12_) );
	DFFPOSX1 DFFPOSX1_1095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_17362__13_), .Q(registers_r31_13_) );
	DFFPOSX1 DFFPOSX1_1096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_17362__14_), .Q(registers_r31_14_) );
	DFFPOSX1 DFFPOSX1_1097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_17362__15_), .Q(registers_r31_15_) );
	DFFPOSX1 DFFPOSX1_1098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_17362__16_), .Q(registers_r31_16_) );
	DFFPOSX1 DFFPOSX1_1099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_17362__17_), .Q(registers_r31_17_) );
	DFFPOSX1 DFFPOSX1_1100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_17362__18_), .Q(registers_r31_18_) );
	DFFPOSX1 DFFPOSX1_1101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_17362__19_), .Q(registers_r31_19_) );
	DFFPOSX1 DFFPOSX1_1102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_17362__20_), .Q(registers_r31_20_) );
	DFFPOSX1 DFFPOSX1_1103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_17362__21_), .Q(registers_r31_21_) );
	DFFPOSX1 DFFPOSX1_1104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_17362__22_), .Q(registers_r31_22_) );
	DFFPOSX1 DFFPOSX1_1105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_17362__23_), .Q(registers_r31_23_) );
	DFFPOSX1 DFFPOSX1_1106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_17362__24_), .Q(registers_r31_24_) );
	DFFPOSX1 DFFPOSX1_1107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_17362__25_), .Q(registers_r31_25_) );
	DFFPOSX1 DFFPOSX1_1108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_17362__26_), .Q(registers_r31_26_) );
	DFFPOSX1 DFFPOSX1_1109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_17362__27_), .Q(registers_r31_27_) );
	DFFPOSX1 DFFPOSX1_1110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_17362__28_), .Q(registers_r31_28_) );
	DFFPOSX1 DFFPOSX1_1111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_17362__29_), .Q(registers_r31_29_) );
	DFFPOSX1 DFFPOSX1_1112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_17362__30_), .Q(registers_r31_30_) );
	DFFPOSX1 DFFPOSX1_1113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_17362__31_), .Q(registers_r31_31_) );
endmodule
